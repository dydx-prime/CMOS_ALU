magic
tech sky130A
timestamp 1767404609
<< nwell >>
rect -120 -1945 -30 -1825
rect 470 -1930 560 -1840
rect -120 -2055 340 -1945
rect 470 -2015 830 -1930
rect 100 -2185 340 -2055
rect 590 -2370 830 -2015
rect 965 -1955 1055 -1835
rect 1530 -1845 1710 -1755
rect 2660 -1815 2840 -1725
rect 1620 -1890 1710 -1845
rect 1620 -1955 1770 -1890
rect 2055 -1930 2145 -1840
rect 2750 -1860 2840 -1815
rect 2750 -1925 2900 -1860
rect 3185 -1910 3275 -1790
rect 3775 -1895 3865 -1805
rect 965 -2065 1425 -1955
rect 1620 -1975 1925 -1955
rect 1185 -2195 1425 -2065
rect 1685 -2195 1925 -1975
rect 2055 -2015 2415 -1930
rect 2750 -1945 3055 -1925
rect 2175 -2370 2415 -2015
rect 2815 -2165 3055 -1945
rect 3185 -2020 3645 -1910
rect 3775 -1980 4135 -1895
rect 3405 -2150 3645 -2020
rect 3895 -2335 4135 -1980
rect 4270 -1920 4360 -1800
rect 4835 -1810 5015 -1720
rect 5965 -1780 6145 -1690
rect 4925 -1855 5015 -1810
rect 4925 -1920 5075 -1855
rect 5360 -1895 5450 -1805
rect 6055 -1825 6145 -1780
rect 6055 -1890 6205 -1825
rect 6490 -1875 6580 -1755
rect 7080 -1860 7170 -1770
rect 4270 -2030 4730 -1920
rect 4925 -1940 5230 -1920
rect 4490 -2160 4730 -2030
rect 4990 -2160 5230 -1940
rect 5360 -1980 5720 -1895
rect 6055 -1910 6360 -1890
rect 5480 -2335 5720 -1980
rect 6120 -2130 6360 -1910
rect 6490 -1985 6950 -1875
rect 7080 -1945 7440 -1860
rect 6710 -2115 6950 -1985
rect 7200 -2300 7440 -1945
rect 7575 -1885 7665 -1765
rect 8140 -1775 8320 -1685
rect 9270 -1745 9450 -1655
rect 8230 -1820 8320 -1775
rect 8230 -1885 8380 -1820
rect 8665 -1860 8755 -1770
rect 9360 -1790 9450 -1745
rect 9360 -1855 9510 -1790
rect 9795 -1840 9885 -1720
rect 10385 -1825 10475 -1735
rect 7575 -1995 8035 -1885
rect 8230 -1905 8535 -1885
rect 7795 -2125 8035 -1995
rect 8295 -2125 8535 -1905
rect 8665 -1945 9025 -1860
rect 9360 -1875 9665 -1855
rect 8785 -2300 9025 -1945
rect 9425 -2095 9665 -1875
rect 9795 -1950 10255 -1840
rect 10385 -1910 10745 -1825
rect 10015 -2080 10255 -1950
rect 10505 -2265 10745 -1910
rect 10880 -1850 10970 -1730
rect 11445 -1740 11625 -1650
rect 12575 -1710 12755 -1620
rect 11535 -1785 11625 -1740
rect 11535 -1850 11685 -1785
rect 11970 -1825 12060 -1735
rect 12665 -1755 12755 -1710
rect 12665 -1820 12815 -1755
rect 10880 -1960 11340 -1850
rect 11535 -1870 11840 -1850
rect 11100 -2090 11340 -1960
rect 11600 -2090 11840 -1870
rect 11970 -1910 12330 -1825
rect 12665 -1840 12970 -1820
rect 12090 -2265 12330 -1910
rect 12730 -2060 12970 -1840
rect 95 -2995 275 -2905
rect 185 -3040 275 -2995
rect 915 -2970 1093 -2880
rect 3400 -2960 3580 -2870
rect 185 -3105 335 -3040
rect 185 -3125 490 -3105
rect 915 -3110 1055 -2970
rect 3490 -3005 3580 -2960
rect 4220 -2935 4398 -2845
rect 6705 -2925 6885 -2835
rect 3490 -3070 3640 -3005
rect 3490 -3090 3795 -3070
rect 4220 -3075 4360 -2935
rect 6795 -2970 6885 -2925
rect 7525 -2900 7703 -2810
rect 10010 -2890 10190 -2800
rect 6795 -3035 6945 -2970
rect 6795 -3055 7100 -3035
rect 7525 -3040 7665 -2900
rect 10100 -2935 10190 -2890
rect 10830 -2865 11008 -2775
rect 10100 -3000 10250 -2935
rect 10100 -3020 10405 -3000
rect 10830 -3005 10970 -2865
rect 250 -3345 490 -3125
rect 3555 -3310 3795 -3090
rect 6860 -3275 7100 -3055
rect 10165 -3240 10405 -3020
rect 13185 -3160 13360 -3070
rect 13615 -3120 13790 -3030
rect 910 -3565 1088 -3475
rect 1620 -3495 1800 -3405
rect 1710 -3540 1800 -3495
rect 2440 -3470 2618 -3380
rect 910 -3705 1050 -3565
rect 1710 -3605 1860 -3540
rect 1710 -3625 2015 -3605
rect 2440 -3610 2580 -3470
rect 4215 -3530 4393 -3440
rect 4925 -3460 5105 -3370
rect 5015 -3505 5105 -3460
rect 5745 -3435 5923 -3345
rect 1775 -3845 2015 -3625
rect 4215 -3670 4355 -3530
rect 5015 -3570 5165 -3505
rect 5015 -3590 5320 -3570
rect 5745 -3575 5885 -3435
rect 7520 -3495 7698 -3405
rect 8230 -3425 8410 -3335
rect 8320 -3470 8410 -3425
rect 9050 -3400 9228 -3310
rect 2700 -3765 2875 -3675
rect 2790 -3895 2875 -3765
rect 5080 -3810 5320 -3590
rect 7520 -3635 7660 -3495
rect 8320 -3535 8470 -3470
rect 8320 -3555 8625 -3535
rect 9050 -3540 9190 -3400
rect 10825 -3460 11003 -3370
rect 11535 -3390 11715 -3300
rect 11625 -3435 11715 -3390
rect 12355 -3365 12533 -3275
rect 13275 -3290 13360 -3160
rect 13705 -3250 13790 -3120
rect 6030 -3730 6205 -3640
rect 6120 -3860 6205 -3730
rect 8385 -3775 8625 -3555
rect 10825 -3600 10965 -3460
rect 11625 -3500 11775 -3435
rect 11625 -3520 11930 -3500
rect 12355 -3505 12495 -3365
rect 9345 -3695 9520 -3605
rect 9435 -3825 9520 -3695
rect 11690 -3740 11930 -3520
rect 13275 -3730 13515 -3290
rect 13705 -3690 13945 -3250
rect 2435 -4065 2613 -3975
rect 45 -4255 225 -4165
rect 135 -4300 225 -4255
rect 865 -4230 1043 -4140
rect 2435 -4205 2575 -4065
rect 135 -4365 285 -4300
rect 135 -4385 440 -4365
rect 865 -4370 1005 -4230
rect 2790 -4335 3030 -3895
rect 5740 -4030 5918 -3940
rect 3350 -4220 3530 -4130
rect 3440 -4265 3530 -4220
rect 4170 -4195 4348 -4105
rect 5740 -4170 5880 -4030
rect 3440 -4330 3590 -4265
rect 3440 -4350 3745 -4330
rect 4170 -4335 4310 -4195
rect 6120 -4300 6360 -3860
rect 9045 -3995 9223 -3905
rect 6655 -4185 6835 -4095
rect 6745 -4230 6835 -4185
rect 7475 -4160 7653 -4070
rect 9045 -4135 9185 -3995
rect 6745 -4295 6895 -4230
rect 6745 -4315 7050 -4295
rect 7475 -4300 7615 -4160
rect 9435 -4265 9675 -3825
rect 12350 -3960 12528 -3870
rect 9960 -4150 10140 -4060
rect 10050 -4195 10140 -4150
rect 10780 -4125 10958 -4035
rect 12350 -4100 12490 -3960
rect 10050 -4260 10200 -4195
rect 10050 -4280 10355 -4260
rect 10780 -4265 10920 -4125
rect 200 -4605 440 -4385
rect 3505 -4570 3745 -4350
rect 6810 -4535 7050 -4315
rect 10115 -4500 10355 -4280
rect 860 -4825 1038 -4735
rect 4165 -4790 4343 -4700
rect 7470 -4755 7648 -4665
rect 10775 -4720 10953 -4630
rect 860 -4965 1000 -4825
rect 4165 -4930 4305 -4790
rect 7470 -4895 7610 -4755
rect 10775 -4860 10915 -4720
rect 9325 -5360 9500 -5270
rect 6220 -5480 6395 -5390
rect 2775 -5585 2950 -5495
rect 2865 -5715 2950 -5585
rect 6310 -5610 6395 -5480
rect 9415 -5490 9500 -5360
rect 2865 -6155 3105 -5715
rect 6310 -6050 6550 -5610
rect 9415 -5930 9655 -5490
<< nmos >>
rect 165 -2665 180 -2465
rect 250 -2665 265 -2465
rect 660 -2675 675 -2575
rect 750 -2675 765 -2575
rect 1255 -2675 1270 -2475
rect 1335 -2675 1350 -2475
rect 1800 -2675 1815 -2575
rect 2245 -2675 2260 -2575
rect 2335 -2675 2350 -2575
rect 2930 -2645 2945 -2545
rect 3470 -2630 3485 -2430
rect 3555 -2630 3570 -2430
rect 3965 -2640 3980 -2540
rect 4055 -2640 4070 -2540
rect 4560 -2640 4575 -2440
rect 4640 -2640 4655 -2440
rect 5105 -2640 5120 -2540
rect 5550 -2640 5565 -2540
rect 5640 -2640 5655 -2540
rect 6235 -2610 6250 -2510
rect 6775 -2595 6790 -2395
rect 6860 -2595 6875 -2395
rect 7270 -2605 7285 -2505
rect 7360 -2605 7375 -2505
rect 7865 -2605 7880 -2405
rect 7945 -2605 7960 -2405
rect 8410 -2605 8425 -2505
rect 8855 -2605 8870 -2505
rect 8945 -2605 8960 -2505
rect 9540 -2575 9555 -2475
rect 10080 -2560 10095 -2360
rect 10165 -2560 10180 -2360
rect 10575 -2570 10590 -2470
rect 10665 -2570 10680 -2470
rect 11170 -2570 11185 -2370
rect 11250 -2570 11265 -2370
rect 11715 -2570 11730 -2470
rect 12160 -2570 12175 -2470
rect 12250 -2570 12265 -2470
rect 12845 -2540 12860 -2440
rect 980 -3290 995 -3190
rect 4285 -3255 4300 -3155
rect 365 -3825 380 -3725
rect 975 -3885 990 -3785
rect 7590 -3220 7605 -3120
rect 2505 -3790 2520 -3690
rect 3670 -3790 3685 -3690
rect 4280 -3850 4295 -3750
rect 1890 -4325 1905 -4225
rect 2500 -4385 2515 -4285
rect 10895 -3185 10910 -3085
rect 5810 -3755 5825 -3655
rect 6975 -3755 6990 -3655
rect 7585 -3815 7600 -3715
rect 5195 -4290 5210 -4190
rect 930 -4550 945 -4450
rect 2900 -4715 2915 -4515
rect 5805 -4350 5820 -4250
rect 9115 -3720 9130 -3620
rect 10280 -3720 10295 -3620
rect 10890 -3780 10905 -3680
rect 8500 -4255 8515 -4155
rect 4235 -4515 4250 -4415
rect 6230 -4680 6245 -4480
rect 9110 -4315 9125 -4215
rect 12420 -3685 12435 -3585
rect 11805 -4220 11820 -4120
rect 13385 -4110 13400 -3910
rect 13815 -4070 13830 -3870
rect 7540 -4480 7555 -4380
rect 9545 -4645 9560 -4445
rect 12415 -4280 12430 -4180
rect 10845 -4445 10860 -4345
rect 315 -5085 330 -4985
rect 925 -5145 940 -5045
rect 3620 -5050 3635 -4950
rect 4230 -5110 4245 -5010
rect 6925 -5015 6940 -4915
rect 7535 -5075 7550 -4975
rect 10230 -4980 10245 -4880
rect 10840 -5040 10855 -4940
rect 2975 -6535 2990 -6335
rect 6420 -6430 6435 -6230
rect 9525 -6310 9540 -6110
<< pmos >>
rect 165 -2165 180 -1965
rect 250 -2165 265 -1965
rect 660 -2350 675 -1950
rect 750 -2350 765 -1950
rect 1255 -2175 1270 -1975
rect 1335 -2175 1350 -1975
rect 1800 -2175 1815 -1975
rect 2245 -2350 2260 -1950
rect 2335 -2350 2350 -1950
rect 2930 -2145 2945 -1945
rect 3470 -2130 3485 -1930
rect 3555 -2130 3570 -1930
rect 3965 -2315 3980 -1915
rect 4055 -2315 4070 -1915
rect 4560 -2140 4575 -1940
rect 4640 -2140 4655 -1940
rect 5105 -2140 5120 -1940
rect 5550 -2315 5565 -1915
rect 5640 -2315 5655 -1915
rect 6235 -2110 6250 -1910
rect 6775 -2095 6790 -1895
rect 6860 -2095 6875 -1895
rect 7270 -2280 7285 -1880
rect 7360 -2280 7375 -1880
rect 7865 -2105 7880 -1905
rect 7945 -2105 7960 -1905
rect 8410 -2105 8425 -1905
rect 8855 -2280 8870 -1880
rect 8945 -2280 8960 -1880
rect 9540 -2075 9555 -1875
rect 10080 -2060 10095 -1860
rect 10165 -2060 10180 -1860
rect 10575 -2245 10590 -1845
rect 10665 -2245 10680 -1845
rect 11170 -2070 11185 -1870
rect 11250 -2070 11265 -1870
rect 11715 -2070 11730 -1870
rect 12160 -2245 12175 -1845
rect 12250 -2245 12265 -1845
rect 12845 -2040 12860 -1840
rect 980 -3090 995 -2990
rect 4285 -3055 4300 -2955
rect 7590 -3020 7605 -2920
rect 10895 -2985 10910 -2885
rect 365 -3325 380 -3125
rect 3670 -3290 3685 -3090
rect 975 -3685 990 -3585
rect 2505 -3590 2520 -3490
rect 6975 -3255 6990 -3055
rect 1890 -3825 1905 -3625
rect 4280 -3650 4295 -3550
rect 5810 -3555 5825 -3455
rect 10280 -3220 10295 -3020
rect 5195 -3790 5210 -3590
rect 2500 -4185 2515 -4085
rect 930 -4350 945 -4250
rect 315 -4585 330 -4385
rect 2900 -4315 2915 -3915
rect 7585 -3615 7600 -3515
rect 9115 -3520 9130 -3420
rect 8500 -3755 8515 -3555
rect 5805 -4150 5820 -4050
rect 4235 -4315 4250 -4215
rect 3620 -4550 3635 -4350
rect 6230 -4280 6245 -3880
rect 10890 -3580 10905 -3480
rect 12420 -3485 12435 -3385
rect 11805 -3720 11820 -3520
rect 9110 -4115 9125 -4015
rect 7540 -4280 7555 -4180
rect 6925 -4515 6940 -4315
rect 9545 -4245 9560 -3845
rect 13385 -3710 13400 -3310
rect 13815 -3670 13830 -3270
rect 12415 -4080 12430 -3980
rect 10845 -4245 10860 -4145
rect 10230 -4480 10245 -4280
rect 925 -4945 940 -4845
rect 4230 -4910 4245 -4810
rect 7535 -4875 7550 -4775
rect 10840 -4840 10855 -4740
rect 2975 -6135 2990 -5735
rect 6420 -6030 6435 -5630
rect 9525 -5910 9540 -5510
<< ndiff >>
rect 120 -2505 165 -2465
rect 120 -2615 125 -2505
rect 150 -2615 165 -2505
rect 120 -2665 165 -2615
rect 180 -2665 250 -2465
rect 265 -2500 320 -2465
rect 265 -2610 290 -2500
rect 315 -2610 320 -2500
rect 1205 -2515 1255 -2475
rect 265 -2665 320 -2610
rect 610 -2595 660 -2575
rect 610 -2655 615 -2595
rect 640 -2655 660 -2595
rect 610 -2675 660 -2655
rect 675 -2595 750 -2575
rect 675 -2655 700 -2595
rect 725 -2655 750 -2595
rect 675 -2675 750 -2655
rect 765 -2595 810 -2575
rect 765 -2655 775 -2595
rect 800 -2655 810 -2595
rect 765 -2675 810 -2655
rect 1205 -2625 1210 -2515
rect 1235 -2625 1255 -2515
rect 1205 -2675 1255 -2625
rect 1270 -2675 1335 -2475
rect 1350 -2510 1405 -2475
rect 1350 -2620 1375 -2510
rect 1400 -2620 1405 -2510
rect 3425 -2470 3470 -2430
rect 2835 -2560 2930 -2545
rect 1350 -2675 1405 -2620
rect 1705 -2590 1800 -2575
rect 1705 -2660 1735 -2590
rect 1765 -2660 1800 -2590
rect 1705 -2675 1800 -2660
rect 1815 -2590 1905 -2575
rect 1815 -2660 1845 -2590
rect 1875 -2660 1905 -2590
rect 1815 -2675 1905 -2660
rect 2195 -2595 2245 -2575
rect 2195 -2655 2200 -2595
rect 2225 -2655 2245 -2595
rect 2195 -2675 2245 -2655
rect 2260 -2595 2335 -2575
rect 2260 -2655 2285 -2595
rect 2310 -2655 2335 -2595
rect 2260 -2675 2335 -2655
rect 2350 -2595 2395 -2575
rect 2350 -2655 2360 -2595
rect 2385 -2655 2395 -2595
rect 2835 -2630 2865 -2560
rect 2895 -2630 2930 -2560
rect 2835 -2645 2930 -2630
rect 2945 -2560 3035 -2545
rect 2945 -2630 2975 -2560
rect 3005 -2630 3035 -2560
rect 3425 -2580 3430 -2470
rect 3455 -2580 3470 -2470
rect 3425 -2630 3470 -2580
rect 3485 -2630 3555 -2430
rect 3570 -2465 3625 -2430
rect 3570 -2575 3595 -2465
rect 3620 -2575 3625 -2465
rect 4510 -2480 4560 -2440
rect 3570 -2630 3625 -2575
rect 3915 -2560 3965 -2540
rect 3915 -2620 3920 -2560
rect 3945 -2620 3965 -2560
rect 2945 -2645 3035 -2630
rect 2350 -2675 2395 -2655
rect 3915 -2640 3965 -2620
rect 3980 -2560 4055 -2540
rect 3980 -2620 4005 -2560
rect 4030 -2620 4055 -2560
rect 3980 -2640 4055 -2620
rect 4070 -2560 4115 -2540
rect 4070 -2620 4080 -2560
rect 4105 -2620 4115 -2560
rect 4070 -2640 4115 -2620
rect 4510 -2590 4515 -2480
rect 4540 -2590 4560 -2480
rect 4510 -2640 4560 -2590
rect 4575 -2640 4640 -2440
rect 4655 -2475 4710 -2440
rect 4655 -2585 4680 -2475
rect 4705 -2585 4710 -2475
rect 6730 -2435 6775 -2395
rect 6140 -2525 6235 -2510
rect 4655 -2640 4710 -2585
rect 5010 -2555 5105 -2540
rect 5010 -2625 5040 -2555
rect 5070 -2625 5105 -2555
rect 5010 -2640 5105 -2625
rect 5120 -2555 5210 -2540
rect 5120 -2625 5150 -2555
rect 5180 -2625 5210 -2555
rect 5120 -2640 5210 -2625
rect 5500 -2560 5550 -2540
rect 5500 -2620 5505 -2560
rect 5530 -2620 5550 -2560
rect 5500 -2640 5550 -2620
rect 5565 -2560 5640 -2540
rect 5565 -2620 5590 -2560
rect 5615 -2620 5640 -2560
rect 5565 -2640 5640 -2620
rect 5655 -2560 5700 -2540
rect 5655 -2620 5665 -2560
rect 5690 -2620 5700 -2560
rect 6140 -2595 6170 -2525
rect 6200 -2595 6235 -2525
rect 6140 -2610 6235 -2595
rect 6250 -2525 6340 -2510
rect 6250 -2595 6280 -2525
rect 6310 -2595 6340 -2525
rect 6730 -2545 6735 -2435
rect 6760 -2545 6775 -2435
rect 6730 -2595 6775 -2545
rect 6790 -2595 6860 -2395
rect 6875 -2430 6930 -2395
rect 6875 -2540 6900 -2430
rect 6925 -2540 6930 -2430
rect 7815 -2445 7865 -2405
rect 6875 -2595 6930 -2540
rect 7220 -2525 7270 -2505
rect 7220 -2585 7225 -2525
rect 7250 -2585 7270 -2525
rect 6250 -2610 6340 -2595
rect 5655 -2640 5700 -2620
rect 7220 -2605 7270 -2585
rect 7285 -2525 7360 -2505
rect 7285 -2585 7310 -2525
rect 7335 -2585 7360 -2525
rect 7285 -2605 7360 -2585
rect 7375 -2525 7420 -2505
rect 7375 -2585 7385 -2525
rect 7410 -2585 7420 -2525
rect 7375 -2605 7420 -2585
rect 7815 -2555 7820 -2445
rect 7845 -2555 7865 -2445
rect 7815 -2605 7865 -2555
rect 7880 -2605 7945 -2405
rect 7960 -2440 8015 -2405
rect 7960 -2550 7985 -2440
rect 8010 -2550 8015 -2440
rect 10035 -2400 10080 -2360
rect 9445 -2490 9540 -2475
rect 7960 -2605 8015 -2550
rect 8315 -2520 8410 -2505
rect 8315 -2590 8345 -2520
rect 8375 -2590 8410 -2520
rect 8315 -2605 8410 -2590
rect 8425 -2520 8515 -2505
rect 8425 -2590 8455 -2520
rect 8485 -2590 8515 -2520
rect 8425 -2605 8515 -2590
rect 8805 -2525 8855 -2505
rect 8805 -2585 8810 -2525
rect 8835 -2585 8855 -2525
rect 8805 -2605 8855 -2585
rect 8870 -2525 8945 -2505
rect 8870 -2585 8895 -2525
rect 8920 -2585 8945 -2525
rect 8870 -2605 8945 -2585
rect 8960 -2525 9005 -2505
rect 8960 -2585 8970 -2525
rect 8995 -2585 9005 -2525
rect 9445 -2560 9475 -2490
rect 9505 -2560 9540 -2490
rect 9445 -2575 9540 -2560
rect 9555 -2490 9645 -2475
rect 9555 -2560 9585 -2490
rect 9615 -2560 9645 -2490
rect 10035 -2510 10040 -2400
rect 10065 -2510 10080 -2400
rect 10035 -2560 10080 -2510
rect 10095 -2560 10165 -2360
rect 10180 -2395 10235 -2360
rect 10180 -2505 10205 -2395
rect 10230 -2505 10235 -2395
rect 11120 -2410 11170 -2370
rect 10180 -2560 10235 -2505
rect 10525 -2490 10575 -2470
rect 10525 -2550 10530 -2490
rect 10555 -2550 10575 -2490
rect 9555 -2575 9645 -2560
rect 8960 -2605 9005 -2585
rect 10525 -2570 10575 -2550
rect 10590 -2490 10665 -2470
rect 10590 -2550 10615 -2490
rect 10640 -2550 10665 -2490
rect 10590 -2570 10665 -2550
rect 10680 -2490 10725 -2470
rect 10680 -2550 10690 -2490
rect 10715 -2550 10725 -2490
rect 10680 -2570 10725 -2550
rect 11120 -2520 11125 -2410
rect 11150 -2520 11170 -2410
rect 11120 -2570 11170 -2520
rect 11185 -2570 11250 -2370
rect 11265 -2405 11320 -2370
rect 11265 -2515 11290 -2405
rect 11315 -2515 11320 -2405
rect 12750 -2455 12845 -2440
rect 11265 -2570 11320 -2515
rect 11620 -2485 11715 -2470
rect 11620 -2555 11650 -2485
rect 11680 -2555 11715 -2485
rect 11620 -2570 11715 -2555
rect 11730 -2485 11820 -2470
rect 11730 -2555 11760 -2485
rect 11790 -2555 11820 -2485
rect 11730 -2570 11820 -2555
rect 12110 -2490 12160 -2470
rect 12110 -2550 12115 -2490
rect 12140 -2550 12160 -2490
rect 12110 -2570 12160 -2550
rect 12175 -2490 12250 -2470
rect 12175 -2550 12200 -2490
rect 12225 -2550 12250 -2490
rect 12175 -2570 12250 -2550
rect 12265 -2490 12310 -2470
rect 12265 -2550 12275 -2490
rect 12300 -2550 12310 -2490
rect 12750 -2525 12780 -2455
rect 12810 -2525 12845 -2455
rect 12750 -2540 12845 -2525
rect 12860 -2455 12950 -2440
rect 12860 -2525 12890 -2455
rect 12920 -2525 12950 -2455
rect 12860 -2540 12950 -2525
rect 12265 -2570 12310 -2550
rect 935 -3200 980 -3190
rect 935 -3280 945 -3200
rect 965 -3280 980 -3200
rect 935 -3290 980 -3280
rect 995 -3200 1035 -3190
rect 995 -3280 1010 -3200
rect 1030 -3280 1035 -3200
rect 995 -3290 1035 -3280
rect 4240 -3165 4285 -3155
rect 4240 -3245 4250 -3165
rect 4270 -3245 4285 -3165
rect 4240 -3255 4285 -3245
rect 4300 -3165 4340 -3155
rect 4300 -3245 4315 -3165
rect 4335 -3245 4340 -3165
rect 4300 -3255 4340 -3245
rect 270 -3740 365 -3725
rect 270 -3810 300 -3740
rect 330 -3810 365 -3740
rect 270 -3825 365 -3810
rect 380 -3740 470 -3725
rect 380 -3810 410 -3740
rect 440 -3810 470 -3740
rect 380 -3825 470 -3810
rect 930 -3795 975 -3785
rect 930 -3875 940 -3795
rect 960 -3875 975 -3795
rect 930 -3885 975 -3875
rect 990 -3795 1030 -3785
rect 990 -3875 1005 -3795
rect 1025 -3875 1030 -3795
rect 990 -3885 1030 -3875
rect 7545 -3130 7590 -3120
rect 7545 -3210 7555 -3130
rect 7575 -3210 7590 -3130
rect 7545 -3220 7590 -3210
rect 7605 -3130 7645 -3120
rect 7605 -3210 7620 -3130
rect 7640 -3210 7645 -3130
rect 7605 -3220 7645 -3210
rect 2460 -3700 2505 -3690
rect 2460 -3780 2470 -3700
rect 2490 -3780 2505 -3700
rect 2460 -3790 2505 -3780
rect 2520 -3700 2560 -3690
rect 2520 -3780 2535 -3700
rect 2555 -3780 2560 -3700
rect 3575 -3705 3670 -3690
rect 2520 -3790 2560 -3780
rect 3575 -3775 3605 -3705
rect 3635 -3775 3670 -3705
rect 3575 -3790 3670 -3775
rect 3685 -3705 3775 -3690
rect 3685 -3775 3715 -3705
rect 3745 -3775 3775 -3705
rect 3685 -3790 3775 -3775
rect 4235 -3760 4280 -3750
rect 4235 -3840 4245 -3760
rect 4265 -3840 4280 -3760
rect 4235 -3850 4280 -3840
rect 4295 -3760 4335 -3750
rect 4295 -3840 4310 -3760
rect 4330 -3840 4335 -3760
rect 4295 -3850 4335 -3840
rect 1795 -4240 1890 -4225
rect 1795 -4310 1825 -4240
rect 1855 -4310 1890 -4240
rect 1795 -4325 1890 -4310
rect 1905 -4240 1995 -4225
rect 1905 -4310 1935 -4240
rect 1965 -4310 1995 -4240
rect 1905 -4325 1995 -4310
rect 2455 -4295 2500 -4285
rect 2455 -4375 2465 -4295
rect 2485 -4375 2500 -4295
rect 2455 -4385 2500 -4375
rect 2515 -4295 2555 -4285
rect 2515 -4375 2530 -4295
rect 2550 -4375 2555 -4295
rect 10850 -3095 10895 -3085
rect 10850 -3175 10860 -3095
rect 10880 -3175 10895 -3095
rect 10850 -3185 10895 -3175
rect 10910 -3095 10950 -3085
rect 10910 -3175 10925 -3095
rect 10945 -3175 10950 -3095
rect 10910 -3185 10950 -3175
rect 5765 -3665 5810 -3655
rect 5765 -3745 5775 -3665
rect 5795 -3745 5810 -3665
rect 5765 -3755 5810 -3745
rect 5825 -3665 5865 -3655
rect 5825 -3745 5840 -3665
rect 5860 -3745 5865 -3665
rect 6880 -3670 6975 -3655
rect 5825 -3755 5865 -3745
rect 6880 -3740 6910 -3670
rect 6940 -3740 6975 -3670
rect 6880 -3755 6975 -3740
rect 6990 -3670 7080 -3655
rect 6990 -3740 7020 -3670
rect 7050 -3740 7080 -3670
rect 6990 -3755 7080 -3740
rect 7540 -3725 7585 -3715
rect 7540 -3805 7550 -3725
rect 7570 -3805 7585 -3725
rect 7540 -3815 7585 -3805
rect 7600 -3725 7640 -3715
rect 7600 -3805 7615 -3725
rect 7635 -3805 7640 -3725
rect 7600 -3815 7640 -3805
rect 5100 -4205 5195 -4190
rect 2515 -4385 2555 -4375
rect 5100 -4275 5130 -4205
rect 5160 -4275 5195 -4205
rect 5100 -4290 5195 -4275
rect 5210 -4205 5300 -4190
rect 5210 -4275 5240 -4205
rect 5270 -4275 5300 -4205
rect 5210 -4290 5300 -4275
rect 5760 -4260 5805 -4250
rect 885 -4460 930 -4450
rect 885 -4540 895 -4460
rect 915 -4540 930 -4460
rect 885 -4550 930 -4540
rect 945 -4460 985 -4450
rect 945 -4540 960 -4460
rect 980 -4540 985 -4460
rect 945 -4550 985 -4540
rect 2810 -4545 2900 -4515
rect 2810 -4700 2820 -4545
rect 2875 -4700 2900 -4545
rect 2810 -4715 2900 -4700
rect 2915 -4545 3010 -4515
rect 2915 -4700 2945 -4545
rect 3000 -4700 3010 -4545
rect 5760 -4340 5770 -4260
rect 5790 -4340 5805 -4260
rect 5760 -4350 5805 -4340
rect 5820 -4260 5860 -4250
rect 5820 -4340 5835 -4260
rect 5855 -4340 5860 -4260
rect 9070 -3630 9115 -3620
rect 9070 -3710 9080 -3630
rect 9100 -3710 9115 -3630
rect 9070 -3720 9115 -3710
rect 9130 -3630 9170 -3620
rect 9130 -3710 9145 -3630
rect 9165 -3710 9170 -3630
rect 10185 -3635 10280 -3620
rect 9130 -3720 9170 -3710
rect 10185 -3705 10215 -3635
rect 10245 -3705 10280 -3635
rect 10185 -3720 10280 -3705
rect 10295 -3635 10385 -3620
rect 10295 -3705 10325 -3635
rect 10355 -3705 10385 -3635
rect 10295 -3720 10385 -3705
rect 10845 -3690 10890 -3680
rect 10845 -3770 10855 -3690
rect 10875 -3770 10890 -3690
rect 10845 -3780 10890 -3770
rect 10905 -3690 10945 -3680
rect 10905 -3770 10920 -3690
rect 10940 -3770 10945 -3690
rect 10905 -3780 10945 -3770
rect 8405 -4170 8500 -4155
rect 5820 -4350 5860 -4340
rect 8405 -4240 8435 -4170
rect 8465 -4240 8500 -4170
rect 8405 -4255 8500 -4240
rect 8515 -4170 8605 -4155
rect 8515 -4240 8545 -4170
rect 8575 -4240 8605 -4170
rect 8515 -4255 8605 -4240
rect 9065 -4225 9110 -4215
rect 2915 -4715 3010 -4700
rect 4190 -4425 4235 -4415
rect 4190 -4505 4200 -4425
rect 4220 -4505 4235 -4425
rect 4190 -4515 4235 -4505
rect 4250 -4425 4290 -4415
rect 4250 -4505 4265 -4425
rect 4285 -4505 4290 -4425
rect 4250 -4515 4290 -4505
rect 6140 -4510 6230 -4480
rect 6140 -4665 6150 -4510
rect 6205 -4665 6230 -4510
rect 6140 -4680 6230 -4665
rect 6245 -4510 6340 -4480
rect 6245 -4665 6275 -4510
rect 6330 -4665 6340 -4510
rect 9065 -4305 9075 -4225
rect 9095 -4305 9110 -4225
rect 9065 -4315 9110 -4305
rect 9125 -4225 9165 -4215
rect 9125 -4305 9140 -4225
rect 9160 -4305 9165 -4225
rect 12375 -3595 12420 -3585
rect 12375 -3675 12385 -3595
rect 12405 -3675 12420 -3595
rect 12375 -3685 12420 -3675
rect 12435 -3595 12475 -3585
rect 12435 -3675 12450 -3595
rect 12470 -3675 12475 -3595
rect 12435 -3685 12475 -3675
rect 13725 -3900 13815 -3870
rect 13295 -3940 13385 -3910
rect 11710 -4135 11805 -4120
rect 9125 -4315 9165 -4305
rect 11710 -4205 11740 -4135
rect 11770 -4205 11805 -4135
rect 11710 -4220 11805 -4205
rect 11820 -4135 11910 -4120
rect 13295 -4095 13305 -3940
rect 13360 -4095 13385 -3940
rect 13295 -4110 13385 -4095
rect 13400 -3940 13495 -3910
rect 13400 -4095 13430 -3940
rect 13485 -4095 13495 -3940
rect 13725 -4055 13735 -3900
rect 13790 -4055 13815 -3900
rect 13725 -4070 13815 -4055
rect 13830 -3900 13925 -3870
rect 13830 -4055 13860 -3900
rect 13915 -4055 13925 -3900
rect 13830 -4070 13925 -4055
rect 13400 -4110 13495 -4095
rect 11820 -4205 11850 -4135
rect 11880 -4205 11910 -4135
rect 11820 -4220 11910 -4205
rect 12370 -4190 12415 -4180
rect 6245 -4680 6340 -4665
rect 7495 -4390 7540 -4380
rect 7495 -4470 7505 -4390
rect 7525 -4470 7540 -4390
rect 7495 -4480 7540 -4470
rect 7555 -4390 7595 -4380
rect 7555 -4470 7570 -4390
rect 7590 -4470 7595 -4390
rect 7555 -4480 7595 -4470
rect 9455 -4475 9545 -4445
rect 9455 -4630 9465 -4475
rect 9520 -4630 9545 -4475
rect 9455 -4645 9545 -4630
rect 9560 -4475 9655 -4445
rect 9560 -4630 9590 -4475
rect 9645 -4630 9655 -4475
rect 12370 -4270 12380 -4190
rect 12400 -4270 12415 -4190
rect 12370 -4280 12415 -4270
rect 12430 -4190 12470 -4180
rect 12430 -4270 12445 -4190
rect 12465 -4270 12470 -4190
rect 12430 -4280 12470 -4270
rect 9560 -4645 9655 -4630
rect 10800 -4355 10845 -4345
rect 10800 -4435 10810 -4355
rect 10830 -4435 10845 -4355
rect 10800 -4445 10845 -4435
rect 10860 -4355 10900 -4345
rect 10860 -4435 10875 -4355
rect 10895 -4435 10900 -4355
rect 10860 -4445 10900 -4435
rect 220 -5000 315 -4985
rect 220 -5070 250 -5000
rect 280 -5070 315 -5000
rect 220 -5085 315 -5070
rect 330 -5000 420 -4985
rect 3525 -4965 3620 -4950
rect 330 -5070 360 -5000
rect 390 -5070 420 -5000
rect 3525 -5035 3555 -4965
rect 3585 -5035 3620 -4965
rect 330 -5085 420 -5070
rect 880 -5055 925 -5045
rect 880 -5135 890 -5055
rect 910 -5135 925 -5055
rect 880 -5145 925 -5135
rect 940 -5055 980 -5045
rect 3525 -5050 3620 -5035
rect 3635 -4965 3725 -4950
rect 6830 -4930 6925 -4915
rect 3635 -5035 3665 -4965
rect 3695 -5035 3725 -4965
rect 6830 -5000 6860 -4930
rect 6890 -5000 6925 -4930
rect 3635 -5050 3725 -5035
rect 4185 -5020 4230 -5010
rect 940 -5135 955 -5055
rect 975 -5135 980 -5055
rect 940 -5145 980 -5135
rect 4185 -5100 4195 -5020
rect 4215 -5100 4230 -5020
rect 4185 -5110 4230 -5100
rect 4245 -5020 4285 -5010
rect 6830 -5015 6925 -5000
rect 6940 -4930 7030 -4915
rect 10135 -4895 10230 -4880
rect 6940 -5000 6970 -4930
rect 7000 -5000 7030 -4930
rect 10135 -4965 10165 -4895
rect 10195 -4965 10230 -4895
rect 6940 -5015 7030 -5000
rect 7490 -4985 7535 -4975
rect 4245 -5100 4260 -5020
rect 4280 -5100 4285 -5020
rect 4245 -5110 4285 -5100
rect 7490 -5065 7500 -4985
rect 7520 -5065 7535 -4985
rect 7490 -5075 7535 -5065
rect 7550 -4985 7590 -4975
rect 10135 -4980 10230 -4965
rect 10245 -4895 10335 -4880
rect 10245 -4965 10275 -4895
rect 10305 -4965 10335 -4895
rect 10245 -4980 10335 -4965
rect 10795 -4950 10840 -4940
rect 7550 -5065 7565 -4985
rect 7585 -5065 7590 -4985
rect 7550 -5075 7590 -5065
rect 10795 -5030 10805 -4950
rect 10825 -5030 10840 -4950
rect 10795 -5040 10840 -5030
rect 10855 -4950 10895 -4940
rect 10855 -5030 10870 -4950
rect 10890 -5030 10895 -4950
rect 10855 -5040 10895 -5030
rect 9435 -6140 9525 -6110
rect 6330 -6260 6420 -6230
rect 2885 -6365 2975 -6335
rect 2885 -6520 2895 -6365
rect 2950 -6520 2975 -6365
rect 2885 -6535 2975 -6520
rect 2990 -6365 3085 -6335
rect 2990 -6520 3020 -6365
rect 3075 -6520 3085 -6365
rect 6330 -6415 6340 -6260
rect 6395 -6415 6420 -6260
rect 6330 -6430 6420 -6415
rect 6435 -6260 6530 -6230
rect 6435 -6415 6465 -6260
rect 6520 -6415 6530 -6260
rect 9435 -6295 9445 -6140
rect 9500 -6295 9525 -6140
rect 9435 -6310 9525 -6295
rect 9540 -6140 9635 -6110
rect 9540 -6295 9570 -6140
rect 9625 -6295 9635 -6140
rect 9540 -6310 9635 -6295
rect 6435 -6430 6530 -6415
rect 2990 -6535 3085 -6520
<< pdiff >>
rect 120 -2010 165 -1965
rect 120 -2120 130 -2010
rect 155 -2120 165 -2010
rect 120 -2165 165 -2120
rect 180 -2010 250 -1965
rect 180 -2120 205 -2010
rect 230 -2120 250 -2010
rect 180 -2165 250 -2120
rect 265 -2010 315 -1965
rect 265 -2120 285 -2010
rect 310 -2120 315 -2010
rect 265 -2165 315 -2120
rect 610 -2020 660 -1950
rect 610 -2220 615 -2020
rect 645 -2220 660 -2020
rect 610 -2350 660 -2220
rect 675 -2350 750 -1950
rect 765 -2015 810 -1950
rect 765 -2215 775 -2015
rect 805 -2215 810 -2015
rect 1205 -2020 1255 -1975
rect 1205 -2130 1215 -2020
rect 1240 -2130 1255 -2020
rect 1205 -2175 1255 -2130
rect 1270 -2020 1335 -1975
rect 1270 -2130 1290 -2020
rect 1315 -2130 1335 -2020
rect 1270 -2175 1335 -2130
rect 1350 -2020 1405 -1975
rect 1350 -2130 1370 -2020
rect 1395 -2130 1405 -2020
rect 1350 -2175 1405 -2130
rect 1705 -2045 1800 -1975
rect 1705 -2115 1730 -2045
rect 1760 -2115 1800 -2045
rect 1705 -2175 1800 -2115
rect 1815 -2045 1905 -1975
rect 1815 -2115 1850 -2045
rect 1880 -2115 1905 -2045
rect 1815 -2175 1905 -2115
rect 2195 -2020 2245 -1950
rect 765 -2350 810 -2215
rect 2195 -2220 2200 -2020
rect 2230 -2220 2245 -2020
rect 2195 -2350 2245 -2220
rect 2260 -2350 2335 -1950
rect 2350 -2015 2395 -1950
rect 2350 -2215 2360 -2015
rect 2390 -2215 2395 -2015
rect 2835 -2015 2930 -1945
rect 2835 -2085 2860 -2015
rect 2890 -2085 2930 -2015
rect 2835 -2145 2930 -2085
rect 2945 -2015 3035 -1945
rect 2945 -2085 2980 -2015
rect 3010 -2085 3035 -2015
rect 2945 -2145 3035 -2085
rect 3425 -1975 3470 -1930
rect 3425 -2085 3435 -1975
rect 3460 -2085 3470 -1975
rect 3425 -2130 3470 -2085
rect 3485 -1975 3555 -1930
rect 3485 -2085 3510 -1975
rect 3535 -2085 3555 -1975
rect 3485 -2130 3555 -2085
rect 3570 -1975 3620 -1930
rect 3570 -2085 3590 -1975
rect 3615 -2085 3620 -1975
rect 3570 -2130 3620 -2085
rect 3915 -1985 3965 -1915
rect 2350 -2350 2395 -2215
rect 3915 -2185 3920 -1985
rect 3950 -2185 3965 -1985
rect 3915 -2315 3965 -2185
rect 3980 -2315 4055 -1915
rect 4070 -1980 4115 -1915
rect 4070 -2180 4080 -1980
rect 4110 -2180 4115 -1980
rect 4510 -1985 4560 -1940
rect 4510 -2095 4520 -1985
rect 4545 -2095 4560 -1985
rect 4510 -2140 4560 -2095
rect 4575 -1985 4640 -1940
rect 4575 -2095 4595 -1985
rect 4620 -2095 4640 -1985
rect 4575 -2140 4640 -2095
rect 4655 -1985 4710 -1940
rect 4655 -2095 4675 -1985
rect 4700 -2095 4710 -1985
rect 4655 -2140 4710 -2095
rect 5010 -2010 5105 -1940
rect 5010 -2080 5035 -2010
rect 5065 -2080 5105 -2010
rect 5010 -2140 5105 -2080
rect 5120 -2010 5210 -1940
rect 5120 -2080 5155 -2010
rect 5185 -2080 5210 -2010
rect 5120 -2140 5210 -2080
rect 5500 -1985 5550 -1915
rect 4070 -2315 4115 -2180
rect 5500 -2185 5505 -1985
rect 5535 -2185 5550 -1985
rect 5500 -2315 5550 -2185
rect 5565 -2315 5640 -1915
rect 5655 -1980 5700 -1915
rect 5655 -2180 5665 -1980
rect 5695 -2180 5700 -1980
rect 6140 -1980 6235 -1910
rect 6140 -2050 6165 -1980
rect 6195 -2050 6235 -1980
rect 6140 -2110 6235 -2050
rect 6250 -1980 6340 -1910
rect 6250 -2050 6285 -1980
rect 6315 -2050 6340 -1980
rect 6250 -2110 6340 -2050
rect 6730 -1940 6775 -1895
rect 6730 -2050 6740 -1940
rect 6765 -2050 6775 -1940
rect 6730 -2095 6775 -2050
rect 6790 -1940 6860 -1895
rect 6790 -2050 6815 -1940
rect 6840 -2050 6860 -1940
rect 6790 -2095 6860 -2050
rect 6875 -1940 6925 -1895
rect 6875 -2050 6895 -1940
rect 6920 -2050 6925 -1940
rect 6875 -2095 6925 -2050
rect 7220 -1950 7270 -1880
rect 5655 -2315 5700 -2180
rect 7220 -2150 7225 -1950
rect 7255 -2150 7270 -1950
rect 7220 -2280 7270 -2150
rect 7285 -2280 7360 -1880
rect 7375 -1945 7420 -1880
rect 7375 -2145 7385 -1945
rect 7415 -2145 7420 -1945
rect 7815 -1950 7865 -1905
rect 7815 -2060 7825 -1950
rect 7850 -2060 7865 -1950
rect 7815 -2105 7865 -2060
rect 7880 -1950 7945 -1905
rect 7880 -2060 7900 -1950
rect 7925 -2060 7945 -1950
rect 7880 -2105 7945 -2060
rect 7960 -1950 8015 -1905
rect 7960 -2060 7980 -1950
rect 8005 -2060 8015 -1950
rect 7960 -2105 8015 -2060
rect 8315 -1975 8410 -1905
rect 8315 -2045 8340 -1975
rect 8370 -2045 8410 -1975
rect 8315 -2105 8410 -2045
rect 8425 -1975 8515 -1905
rect 8425 -2045 8460 -1975
rect 8490 -2045 8515 -1975
rect 8425 -2105 8515 -2045
rect 8805 -1950 8855 -1880
rect 7375 -2280 7420 -2145
rect 8805 -2150 8810 -1950
rect 8840 -2150 8855 -1950
rect 8805 -2280 8855 -2150
rect 8870 -2280 8945 -1880
rect 8960 -1945 9005 -1880
rect 8960 -2145 8970 -1945
rect 9000 -2145 9005 -1945
rect 9445 -1945 9540 -1875
rect 9445 -2015 9470 -1945
rect 9500 -2015 9540 -1945
rect 9445 -2075 9540 -2015
rect 9555 -1945 9645 -1875
rect 9555 -2015 9590 -1945
rect 9620 -2015 9645 -1945
rect 9555 -2075 9645 -2015
rect 10035 -1905 10080 -1860
rect 10035 -2015 10045 -1905
rect 10070 -2015 10080 -1905
rect 10035 -2060 10080 -2015
rect 10095 -1905 10165 -1860
rect 10095 -2015 10120 -1905
rect 10145 -2015 10165 -1905
rect 10095 -2060 10165 -2015
rect 10180 -1905 10230 -1860
rect 10180 -2015 10200 -1905
rect 10225 -2015 10230 -1905
rect 10180 -2060 10230 -2015
rect 10525 -1915 10575 -1845
rect 8960 -2280 9005 -2145
rect 10525 -2115 10530 -1915
rect 10560 -2115 10575 -1915
rect 10525 -2245 10575 -2115
rect 10590 -2245 10665 -1845
rect 10680 -1910 10725 -1845
rect 10680 -2110 10690 -1910
rect 10720 -2110 10725 -1910
rect 11120 -1915 11170 -1870
rect 11120 -2025 11130 -1915
rect 11155 -2025 11170 -1915
rect 11120 -2070 11170 -2025
rect 11185 -1915 11250 -1870
rect 11185 -2025 11205 -1915
rect 11230 -2025 11250 -1915
rect 11185 -2070 11250 -2025
rect 11265 -1915 11320 -1870
rect 11265 -2025 11285 -1915
rect 11310 -2025 11320 -1915
rect 11265 -2070 11320 -2025
rect 11620 -1940 11715 -1870
rect 11620 -2010 11645 -1940
rect 11675 -2010 11715 -1940
rect 11620 -2070 11715 -2010
rect 11730 -1940 11820 -1870
rect 11730 -2010 11765 -1940
rect 11795 -2010 11820 -1940
rect 11730 -2070 11820 -2010
rect 12110 -1915 12160 -1845
rect 10680 -2245 10725 -2110
rect 12110 -2115 12115 -1915
rect 12145 -2115 12160 -1915
rect 12110 -2245 12160 -2115
rect 12175 -2245 12250 -1845
rect 12265 -1910 12310 -1845
rect 12265 -2110 12275 -1910
rect 12305 -2110 12310 -1910
rect 12750 -1910 12845 -1840
rect 12750 -1980 12775 -1910
rect 12805 -1980 12845 -1910
rect 12750 -2040 12845 -1980
rect 12860 -1910 12950 -1840
rect 12860 -1980 12895 -1910
rect 12925 -1980 12950 -1910
rect 12860 -2040 12950 -1980
rect 12265 -2245 12310 -2110
rect 10850 -2895 10895 -2885
rect 7545 -2930 7590 -2920
rect 4240 -2965 4285 -2955
rect 935 -3000 980 -2990
rect 935 -3080 945 -3000
rect 965 -3080 980 -3000
rect 935 -3090 980 -3080
rect 995 -3000 1035 -2990
rect 995 -3080 1005 -3000
rect 1025 -3080 1035 -3000
rect 4240 -3045 4250 -2965
rect 4270 -3045 4285 -2965
rect 995 -3090 1035 -3080
rect 4240 -3055 4285 -3045
rect 4300 -2965 4340 -2955
rect 4300 -3045 4310 -2965
rect 4330 -3045 4340 -2965
rect 7545 -3010 7555 -2930
rect 7575 -3010 7590 -2930
rect 4300 -3055 4340 -3045
rect 7545 -3020 7590 -3010
rect 7605 -2930 7645 -2920
rect 7605 -3010 7615 -2930
rect 7635 -3010 7645 -2930
rect 10850 -2975 10860 -2895
rect 10880 -2975 10895 -2895
rect 7605 -3020 7645 -3010
rect 10850 -2985 10895 -2975
rect 10910 -2895 10950 -2885
rect 10910 -2975 10920 -2895
rect 10940 -2975 10950 -2895
rect 10910 -2985 10950 -2975
rect 270 -3195 365 -3125
rect 270 -3265 295 -3195
rect 325 -3265 365 -3195
rect 270 -3325 365 -3265
rect 380 -3195 470 -3125
rect 3575 -3160 3670 -3090
rect 380 -3265 415 -3195
rect 445 -3265 470 -3195
rect 380 -3325 470 -3265
rect 3575 -3230 3600 -3160
rect 3630 -3230 3670 -3160
rect 3575 -3290 3670 -3230
rect 3685 -3160 3775 -3090
rect 6880 -3125 6975 -3055
rect 3685 -3230 3720 -3160
rect 3750 -3230 3775 -3160
rect 3685 -3290 3775 -3230
rect 2460 -3500 2505 -3490
rect 2460 -3580 2470 -3500
rect 2490 -3580 2505 -3500
rect 930 -3595 975 -3585
rect 930 -3675 940 -3595
rect 960 -3675 975 -3595
rect 930 -3685 975 -3675
rect 990 -3595 1030 -3585
rect 990 -3675 1000 -3595
rect 1020 -3675 1030 -3595
rect 2460 -3590 2505 -3580
rect 2520 -3500 2560 -3490
rect 2520 -3580 2530 -3500
rect 2550 -3580 2560 -3500
rect 6880 -3195 6905 -3125
rect 6935 -3195 6975 -3125
rect 6880 -3255 6975 -3195
rect 6990 -3125 7080 -3055
rect 10185 -3090 10280 -3020
rect 6990 -3195 7025 -3125
rect 7055 -3195 7080 -3125
rect 6990 -3255 7080 -3195
rect 5765 -3465 5810 -3455
rect 2520 -3590 2560 -3580
rect 990 -3685 1030 -3675
rect 1795 -3695 1890 -3625
rect 1795 -3765 1820 -3695
rect 1850 -3765 1890 -3695
rect 1795 -3825 1890 -3765
rect 1905 -3695 1995 -3625
rect 1905 -3765 1940 -3695
rect 1970 -3765 1995 -3695
rect 1905 -3825 1995 -3765
rect 5765 -3545 5775 -3465
rect 5795 -3545 5810 -3465
rect 4235 -3560 4280 -3550
rect 4235 -3640 4245 -3560
rect 4265 -3640 4280 -3560
rect 4235 -3650 4280 -3640
rect 4295 -3560 4335 -3550
rect 4295 -3640 4305 -3560
rect 4325 -3640 4335 -3560
rect 5765 -3555 5810 -3545
rect 5825 -3465 5865 -3455
rect 5825 -3545 5835 -3465
rect 5855 -3545 5865 -3465
rect 10185 -3160 10210 -3090
rect 10240 -3160 10280 -3090
rect 10185 -3220 10280 -3160
rect 10295 -3090 10385 -3020
rect 10295 -3160 10330 -3090
rect 10360 -3160 10385 -3090
rect 10295 -3220 10385 -3160
rect 9070 -3430 9115 -3420
rect 5825 -3555 5865 -3545
rect 4295 -3650 4335 -3640
rect 5100 -3660 5195 -3590
rect 5100 -3730 5125 -3660
rect 5155 -3730 5195 -3660
rect 5100 -3790 5195 -3730
rect 5210 -3660 5300 -3590
rect 5210 -3730 5245 -3660
rect 5275 -3730 5300 -3660
rect 5210 -3790 5300 -3730
rect 2810 -3945 2900 -3915
rect 2455 -4095 2500 -4085
rect 2455 -4175 2465 -4095
rect 2485 -4175 2500 -4095
rect 2455 -4185 2500 -4175
rect 2515 -4095 2555 -4085
rect 2515 -4175 2525 -4095
rect 2545 -4175 2555 -4095
rect 2515 -4185 2555 -4175
rect 885 -4260 930 -4250
rect 885 -4340 895 -4260
rect 915 -4340 930 -4260
rect 885 -4350 930 -4340
rect 945 -4260 985 -4250
rect 945 -4340 955 -4260
rect 975 -4340 985 -4260
rect 945 -4350 985 -4340
rect 220 -4455 315 -4385
rect 220 -4525 245 -4455
rect 275 -4525 315 -4455
rect 220 -4585 315 -4525
rect 330 -4455 420 -4385
rect 330 -4525 365 -4455
rect 395 -4525 420 -4455
rect 330 -4585 420 -4525
rect 2810 -4290 2820 -3945
rect 2885 -4290 2900 -3945
rect 2810 -4315 2900 -4290
rect 2915 -3945 3010 -3915
rect 2915 -4290 2935 -3945
rect 3000 -4290 3010 -3945
rect 9070 -3510 9080 -3430
rect 9100 -3510 9115 -3430
rect 7540 -3525 7585 -3515
rect 7540 -3605 7550 -3525
rect 7570 -3605 7585 -3525
rect 7540 -3615 7585 -3605
rect 7600 -3525 7640 -3515
rect 7600 -3605 7610 -3525
rect 7630 -3605 7640 -3525
rect 9070 -3520 9115 -3510
rect 9130 -3430 9170 -3420
rect 9130 -3510 9140 -3430
rect 9160 -3510 9170 -3430
rect 13725 -3300 13815 -3270
rect 13295 -3340 13385 -3310
rect 12375 -3395 12420 -3385
rect 9130 -3520 9170 -3510
rect 7600 -3615 7640 -3605
rect 8405 -3625 8500 -3555
rect 8405 -3695 8430 -3625
rect 8460 -3695 8500 -3625
rect 8405 -3755 8500 -3695
rect 8515 -3625 8605 -3555
rect 8515 -3695 8550 -3625
rect 8580 -3695 8605 -3625
rect 8515 -3755 8605 -3695
rect 6140 -3910 6230 -3880
rect 5760 -4060 5805 -4050
rect 5760 -4140 5770 -4060
rect 5790 -4140 5805 -4060
rect 5760 -4150 5805 -4140
rect 5820 -4060 5860 -4050
rect 5820 -4140 5830 -4060
rect 5850 -4140 5860 -4060
rect 5820 -4150 5860 -4140
rect 2915 -4315 3010 -4290
rect 4190 -4225 4235 -4215
rect 4190 -4305 4200 -4225
rect 4220 -4305 4235 -4225
rect 4190 -4315 4235 -4305
rect 4250 -4225 4290 -4215
rect 4250 -4305 4260 -4225
rect 4280 -4305 4290 -4225
rect 4250 -4315 4290 -4305
rect 3525 -4420 3620 -4350
rect 3525 -4490 3550 -4420
rect 3580 -4490 3620 -4420
rect 3525 -4550 3620 -4490
rect 3635 -4420 3725 -4350
rect 3635 -4490 3670 -4420
rect 3700 -4490 3725 -4420
rect 3635 -4550 3725 -4490
rect 6140 -4255 6150 -3910
rect 6215 -4255 6230 -3910
rect 6140 -4280 6230 -4255
rect 6245 -3910 6340 -3880
rect 6245 -4255 6265 -3910
rect 6330 -4255 6340 -3910
rect 12375 -3475 12385 -3395
rect 12405 -3475 12420 -3395
rect 10845 -3490 10890 -3480
rect 10845 -3570 10855 -3490
rect 10875 -3570 10890 -3490
rect 10845 -3580 10890 -3570
rect 10905 -3490 10945 -3480
rect 10905 -3570 10915 -3490
rect 10935 -3570 10945 -3490
rect 12375 -3485 12420 -3475
rect 12435 -3395 12475 -3385
rect 12435 -3475 12445 -3395
rect 12465 -3475 12475 -3395
rect 12435 -3485 12475 -3475
rect 10905 -3580 10945 -3570
rect 11710 -3590 11805 -3520
rect 11710 -3660 11735 -3590
rect 11765 -3660 11805 -3590
rect 11710 -3720 11805 -3660
rect 11820 -3590 11910 -3520
rect 11820 -3660 11855 -3590
rect 11885 -3660 11910 -3590
rect 11820 -3720 11910 -3660
rect 9455 -3875 9545 -3845
rect 9065 -4025 9110 -4015
rect 9065 -4105 9075 -4025
rect 9095 -4105 9110 -4025
rect 9065 -4115 9110 -4105
rect 9125 -4025 9165 -4015
rect 9125 -4105 9135 -4025
rect 9155 -4105 9165 -4025
rect 9125 -4115 9165 -4105
rect 6245 -4280 6340 -4255
rect 7495 -4190 7540 -4180
rect 7495 -4270 7505 -4190
rect 7525 -4270 7540 -4190
rect 7495 -4280 7540 -4270
rect 7555 -4190 7595 -4180
rect 7555 -4270 7565 -4190
rect 7585 -4270 7595 -4190
rect 7555 -4280 7595 -4270
rect 6830 -4385 6925 -4315
rect 6830 -4455 6855 -4385
rect 6885 -4455 6925 -4385
rect 6830 -4515 6925 -4455
rect 6940 -4385 7030 -4315
rect 6940 -4455 6975 -4385
rect 7005 -4455 7030 -4385
rect 6940 -4515 7030 -4455
rect 9455 -4220 9465 -3875
rect 9530 -4220 9545 -3875
rect 9455 -4245 9545 -4220
rect 9560 -3875 9655 -3845
rect 9560 -4220 9580 -3875
rect 9645 -4220 9655 -3875
rect 13295 -3685 13305 -3340
rect 13370 -3685 13385 -3340
rect 13295 -3710 13385 -3685
rect 13400 -3340 13495 -3310
rect 13400 -3685 13420 -3340
rect 13485 -3685 13495 -3340
rect 13725 -3645 13735 -3300
rect 13800 -3645 13815 -3300
rect 13725 -3670 13815 -3645
rect 13830 -3300 13925 -3270
rect 13830 -3645 13850 -3300
rect 13915 -3645 13925 -3300
rect 13830 -3670 13925 -3645
rect 13400 -3710 13495 -3685
rect 12370 -3990 12415 -3980
rect 12370 -4070 12380 -3990
rect 12400 -4070 12415 -3990
rect 12370 -4080 12415 -4070
rect 12430 -3990 12470 -3980
rect 12430 -4070 12440 -3990
rect 12460 -4070 12470 -3990
rect 12430 -4080 12470 -4070
rect 9560 -4245 9655 -4220
rect 10800 -4155 10845 -4145
rect 10800 -4235 10810 -4155
rect 10830 -4235 10845 -4155
rect 10800 -4245 10845 -4235
rect 10860 -4155 10900 -4145
rect 10860 -4235 10870 -4155
rect 10890 -4235 10900 -4155
rect 10860 -4245 10900 -4235
rect 10135 -4350 10230 -4280
rect 10135 -4420 10160 -4350
rect 10190 -4420 10230 -4350
rect 10135 -4480 10230 -4420
rect 10245 -4350 10335 -4280
rect 10245 -4420 10280 -4350
rect 10310 -4420 10335 -4350
rect 10245 -4480 10335 -4420
rect 880 -4855 925 -4845
rect 880 -4935 890 -4855
rect 910 -4935 925 -4855
rect 880 -4945 925 -4935
rect 940 -4855 980 -4845
rect 940 -4935 950 -4855
rect 970 -4935 980 -4855
rect 940 -4945 980 -4935
rect 4185 -4820 4230 -4810
rect 4185 -4900 4195 -4820
rect 4215 -4900 4230 -4820
rect 4185 -4910 4230 -4900
rect 4245 -4820 4285 -4810
rect 4245 -4900 4255 -4820
rect 4275 -4900 4285 -4820
rect 4245 -4910 4285 -4900
rect 7490 -4785 7535 -4775
rect 7490 -4865 7500 -4785
rect 7520 -4865 7535 -4785
rect 7490 -4875 7535 -4865
rect 7550 -4785 7590 -4775
rect 7550 -4865 7560 -4785
rect 7580 -4865 7590 -4785
rect 7550 -4875 7590 -4865
rect 10795 -4750 10840 -4740
rect 10795 -4830 10805 -4750
rect 10825 -4830 10840 -4750
rect 10795 -4840 10840 -4830
rect 10855 -4750 10895 -4740
rect 10855 -4830 10865 -4750
rect 10885 -4830 10895 -4750
rect 10855 -4840 10895 -4830
rect 9435 -5540 9525 -5510
rect 6330 -5660 6420 -5630
rect 2885 -5765 2975 -5735
rect 2885 -6110 2895 -5765
rect 2960 -6110 2975 -5765
rect 2885 -6135 2975 -6110
rect 2990 -5765 3085 -5735
rect 2990 -6110 3010 -5765
rect 3075 -6110 3085 -5765
rect 6330 -6005 6340 -5660
rect 6405 -6005 6420 -5660
rect 6330 -6030 6420 -6005
rect 6435 -5660 6530 -5630
rect 6435 -6005 6455 -5660
rect 6520 -6005 6530 -5660
rect 9435 -5885 9445 -5540
rect 9510 -5885 9525 -5540
rect 9435 -5910 9525 -5885
rect 9540 -5540 9635 -5510
rect 9540 -5885 9560 -5540
rect 9625 -5885 9635 -5540
rect 9540 -5910 9635 -5885
rect 6435 -6030 6530 -6005
rect 2990 -6135 3085 -6110
<< ndiffc >>
rect 125 -2615 150 -2505
rect 290 -2610 315 -2500
rect 615 -2655 640 -2595
rect 700 -2655 725 -2595
rect 775 -2655 800 -2595
rect 1210 -2625 1235 -2515
rect 1375 -2620 1400 -2510
rect 1735 -2660 1765 -2590
rect 1845 -2660 1875 -2590
rect 2200 -2655 2225 -2595
rect 2285 -2655 2310 -2595
rect 2360 -2655 2385 -2595
rect 2865 -2630 2895 -2560
rect 2975 -2630 3005 -2560
rect 3430 -2580 3455 -2470
rect 3595 -2575 3620 -2465
rect 3920 -2620 3945 -2560
rect 4005 -2620 4030 -2560
rect 4080 -2620 4105 -2560
rect 4515 -2590 4540 -2480
rect 4680 -2585 4705 -2475
rect 5040 -2625 5070 -2555
rect 5150 -2625 5180 -2555
rect 5505 -2620 5530 -2560
rect 5590 -2620 5615 -2560
rect 5665 -2620 5690 -2560
rect 6170 -2595 6200 -2525
rect 6280 -2595 6310 -2525
rect 6735 -2545 6760 -2435
rect 6900 -2540 6925 -2430
rect 7225 -2585 7250 -2525
rect 7310 -2585 7335 -2525
rect 7385 -2585 7410 -2525
rect 7820 -2555 7845 -2445
rect 7985 -2550 8010 -2440
rect 8345 -2590 8375 -2520
rect 8455 -2590 8485 -2520
rect 8810 -2585 8835 -2525
rect 8895 -2585 8920 -2525
rect 8970 -2585 8995 -2525
rect 9475 -2560 9505 -2490
rect 9585 -2560 9615 -2490
rect 10040 -2510 10065 -2400
rect 10205 -2505 10230 -2395
rect 10530 -2550 10555 -2490
rect 10615 -2550 10640 -2490
rect 10690 -2550 10715 -2490
rect 11125 -2520 11150 -2410
rect 11290 -2515 11315 -2405
rect 11650 -2555 11680 -2485
rect 11760 -2555 11790 -2485
rect 12115 -2550 12140 -2490
rect 12200 -2550 12225 -2490
rect 12275 -2550 12300 -2490
rect 12780 -2525 12810 -2455
rect 12890 -2525 12920 -2455
rect 945 -3280 965 -3200
rect 1010 -3280 1030 -3200
rect 4250 -3245 4270 -3165
rect 4315 -3245 4335 -3165
rect 300 -3810 330 -3740
rect 410 -3810 440 -3740
rect 940 -3875 960 -3795
rect 1005 -3875 1025 -3795
rect 7555 -3210 7575 -3130
rect 7620 -3210 7640 -3130
rect 2470 -3780 2490 -3700
rect 2535 -3780 2555 -3700
rect 3605 -3775 3635 -3705
rect 3715 -3775 3745 -3705
rect 4245 -3840 4265 -3760
rect 4310 -3840 4330 -3760
rect 1825 -4310 1855 -4240
rect 1935 -4310 1965 -4240
rect 2465 -4375 2485 -4295
rect 2530 -4375 2550 -4295
rect 10860 -3175 10880 -3095
rect 10925 -3175 10945 -3095
rect 5775 -3745 5795 -3665
rect 5840 -3745 5860 -3665
rect 6910 -3740 6940 -3670
rect 7020 -3740 7050 -3670
rect 7550 -3805 7570 -3725
rect 7615 -3805 7635 -3725
rect 5130 -4275 5160 -4205
rect 5240 -4275 5270 -4205
rect 895 -4540 915 -4460
rect 960 -4540 980 -4460
rect 2820 -4700 2875 -4545
rect 2945 -4700 3000 -4545
rect 5770 -4340 5790 -4260
rect 5835 -4340 5855 -4260
rect 9080 -3710 9100 -3630
rect 9145 -3710 9165 -3630
rect 10215 -3705 10245 -3635
rect 10325 -3705 10355 -3635
rect 10855 -3770 10875 -3690
rect 10920 -3770 10940 -3690
rect 8435 -4240 8465 -4170
rect 8545 -4240 8575 -4170
rect 4200 -4505 4220 -4425
rect 4265 -4505 4285 -4425
rect 6150 -4665 6205 -4510
rect 6275 -4665 6330 -4510
rect 9075 -4305 9095 -4225
rect 9140 -4305 9160 -4225
rect 12385 -3675 12405 -3595
rect 12450 -3675 12470 -3595
rect 11740 -4205 11770 -4135
rect 13305 -4095 13360 -3940
rect 13430 -4095 13485 -3940
rect 13735 -4055 13790 -3900
rect 13860 -4055 13915 -3900
rect 11850 -4205 11880 -4135
rect 7505 -4470 7525 -4390
rect 7570 -4470 7590 -4390
rect 9465 -4630 9520 -4475
rect 9590 -4630 9645 -4475
rect 12380 -4270 12400 -4190
rect 12445 -4270 12465 -4190
rect 10810 -4435 10830 -4355
rect 10875 -4435 10895 -4355
rect 250 -5070 280 -5000
rect 360 -5070 390 -5000
rect 3555 -5035 3585 -4965
rect 890 -5135 910 -5055
rect 3665 -5035 3695 -4965
rect 6860 -5000 6890 -4930
rect 955 -5135 975 -5055
rect 4195 -5100 4215 -5020
rect 6970 -5000 7000 -4930
rect 10165 -4965 10195 -4895
rect 4260 -5100 4280 -5020
rect 7500 -5065 7520 -4985
rect 10275 -4965 10305 -4895
rect 7565 -5065 7585 -4985
rect 10805 -5030 10825 -4950
rect 10870 -5030 10890 -4950
rect 2895 -6520 2950 -6365
rect 3020 -6520 3075 -6365
rect 6340 -6415 6395 -6260
rect 6465 -6415 6520 -6260
rect 9445 -6295 9500 -6140
rect 9570 -6295 9625 -6140
<< pdiffc >>
rect 130 -2120 155 -2010
rect 205 -2120 230 -2010
rect 285 -2120 310 -2010
rect 615 -2220 645 -2020
rect 775 -2215 805 -2015
rect 1215 -2130 1240 -2020
rect 1290 -2130 1315 -2020
rect 1370 -2130 1395 -2020
rect 1730 -2115 1760 -2045
rect 1850 -2115 1880 -2045
rect 2200 -2220 2230 -2020
rect 2360 -2215 2390 -2015
rect 2860 -2085 2890 -2015
rect 2980 -2085 3010 -2015
rect 3435 -2085 3460 -1975
rect 3510 -2085 3535 -1975
rect 3590 -2085 3615 -1975
rect 3920 -2185 3950 -1985
rect 4080 -2180 4110 -1980
rect 4520 -2095 4545 -1985
rect 4595 -2095 4620 -1985
rect 4675 -2095 4700 -1985
rect 5035 -2080 5065 -2010
rect 5155 -2080 5185 -2010
rect 5505 -2185 5535 -1985
rect 5665 -2180 5695 -1980
rect 6165 -2050 6195 -1980
rect 6285 -2050 6315 -1980
rect 6740 -2050 6765 -1940
rect 6815 -2050 6840 -1940
rect 6895 -2050 6920 -1940
rect 7225 -2150 7255 -1950
rect 7385 -2145 7415 -1945
rect 7825 -2060 7850 -1950
rect 7900 -2060 7925 -1950
rect 7980 -2060 8005 -1950
rect 8340 -2045 8370 -1975
rect 8460 -2045 8490 -1975
rect 8810 -2150 8840 -1950
rect 8970 -2145 9000 -1945
rect 9470 -2015 9500 -1945
rect 9590 -2015 9620 -1945
rect 10045 -2015 10070 -1905
rect 10120 -2015 10145 -1905
rect 10200 -2015 10225 -1905
rect 10530 -2115 10560 -1915
rect 10690 -2110 10720 -1910
rect 11130 -2025 11155 -1915
rect 11205 -2025 11230 -1915
rect 11285 -2025 11310 -1915
rect 11645 -2010 11675 -1940
rect 11765 -2010 11795 -1940
rect 12115 -2115 12145 -1915
rect 12275 -2110 12305 -1910
rect 12775 -1980 12805 -1910
rect 12895 -1980 12925 -1910
rect 945 -3080 965 -3000
rect 1005 -3080 1025 -3000
rect 4250 -3045 4270 -2965
rect 4310 -3045 4330 -2965
rect 7555 -3010 7575 -2930
rect 7615 -3010 7635 -2930
rect 10860 -2975 10880 -2895
rect 10920 -2975 10940 -2895
rect 295 -3265 325 -3195
rect 415 -3265 445 -3195
rect 3600 -3230 3630 -3160
rect 3720 -3230 3750 -3160
rect 2470 -3580 2490 -3500
rect 940 -3675 960 -3595
rect 1000 -3675 1020 -3595
rect 2530 -3580 2550 -3500
rect 6905 -3195 6935 -3125
rect 7025 -3195 7055 -3125
rect 1820 -3765 1850 -3695
rect 1940 -3765 1970 -3695
rect 5775 -3545 5795 -3465
rect 4245 -3640 4265 -3560
rect 4305 -3640 4325 -3560
rect 5835 -3545 5855 -3465
rect 10210 -3160 10240 -3090
rect 10330 -3160 10360 -3090
rect 5125 -3730 5155 -3660
rect 5245 -3730 5275 -3660
rect 2465 -4175 2485 -4095
rect 2525 -4175 2545 -4095
rect 895 -4340 915 -4260
rect 955 -4340 975 -4260
rect 245 -4525 275 -4455
rect 365 -4525 395 -4455
rect 2820 -4290 2885 -3945
rect 2935 -4290 3000 -3945
rect 9080 -3510 9100 -3430
rect 7550 -3605 7570 -3525
rect 7610 -3605 7630 -3525
rect 9140 -3510 9160 -3430
rect 8430 -3695 8460 -3625
rect 8550 -3695 8580 -3625
rect 5770 -4140 5790 -4060
rect 5830 -4140 5850 -4060
rect 4200 -4305 4220 -4225
rect 4260 -4305 4280 -4225
rect 3550 -4490 3580 -4420
rect 3670 -4490 3700 -4420
rect 6150 -4255 6215 -3910
rect 6265 -4255 6330 -3910
rect 12385 -3475 12405 -3395
rect 10855 -3570 10875 -3490
rect 10915 -3570 10935 -3490
rect 12445 -3475 12465 -3395
rect 11735 -3660 11765 -3590
rect 11855 -3660 11885 -3590
rect 9075 -4105 9095 -4025
rect 9135 -4105 9155 -4025
rect 7505 -4270 7525 -4190
rect 7565 -4270 7585 -4190
rect 6855 -4455 6885 -4385
rect 6975 -4455 7005 -4385
rect 9465 -4220 9530 -3875
rect 9580 -4220 9645 -3875
rect 13305 -3685 13370 -3340
rect 13420 -3685 13485 -3340
rect 13735 -3645 13800 -3300
rect 13850 -3645 13915 -3300
rect 12380 -4070 12400 -3990
rect 12440 -4070 12460 -3990
rect 10810 -4235 10830 -4155
rect 10870 -4235 10890 -4155
rect 10160 -4420 10190 -4350
rect 10280 -4420 10310 -4350
rect 890 -4935 910 -4855
rect 950 -4935 970 -4855
rect 4195 -4900 4215 -4820
rect 4255 -4900 4275 -4820
rect 7500 -4865 7520 -4785
rect 7560 -4865 7580 -4785
rect 10805 -4830 10825 -4750
rect 10865 -4830 10885 -4750
rect 2895 -6110 2960 -5765
rect 3010 -6110 3075 -5765
rect 6340 -6005 6405 -5660
rect 6455 -6005 6520 -5660
rect 9445 -5885 9510 -5540
rect 9560 -5885 9625 -5540
<< psubdiff >>
rect 10390 -2605 10465 -2590
rect 9855 -2625 9905 -2615
rect 7085 -2640 7160 -2625
rect 6550 -2660 6600 -2650
rect 3780 -2675 3855 -2660
rect 3245 -2695 3295 -2685
rect 475 -2710 550 -2695
rect -60 -2730 -10 -2720
rect -60 -2755 -45 -2730
rect -25 -2755 -10 -2730
rect 475 -2740 490 -2710
rect 535 -2740 550 -2710
rect 2060 -2710 2135 -2695
rect 475 -2755 550 -2740
rect 1025 -2740 1075 -2730
rect -60 -2765 -10 -2755
rect 1025 -2765 1040 -2740
rect 1060 -2765 1075 -2740
rect 1025 -2775 1075 -2765
rect 1565 -2740 1615 -2730
rect 1565 -2765 1580 -2740
rect 1600 -2765 1615 -2740
rect 2060 -2740 2075 -2710
rect 2120 -2740 2135 -2710
rect 2060 -2755 2135 -2740
rect 2695 -2710 2745 -2700
rect 2695 -2735 2710 -2710
rect 2730 -2735 2745 -2710
rect 3245 -2720 3260 -2695
rect 3280 -2720 3295 -2695
rect 3780 -2705 3795 -2675
rect 3840 -2705 3855 -2675
rect 5365 -2675 5440 -2660
rect 3780 -2720 3855 -2705
rect 4330 -2705 4380 -2695
rect 3245 -2730 3295 -2720
rect 4330 -2730 4345 -2705
rect 4365 -2730 4380 -2705
rect 2695 -2745 2745 -2735
rect 4330 -2740 4380 -2730
rect 4870 -2705 4920 -2695
rect 4870 -2730 4885 -2705
rect 4905 -2730 4920 -2705
rect 5365 -2705 5380 -2675
rect 5425 -2705 5440 -2675
rect 5365 -2720 5440 -2705
rect 6000 -2675 6050 -2665
rect 6000 -2700 6015 -2675
rect 6035 -2700 6050 -2675
rect 6550 -2685 6565 -2660
rect 6585 -2685 6600 -2660
rect 7085 -2670 7100 -2640
rect 7145 -2670 7160 -2640
rect 8670 -2640 8745 -2625
rect 7085 -2685 7160 -2670
rect 7635 -2670 7685 -2660
rect 6550 -2695 6600 -2685
rect 7635 -2695 7650 -2670
rect 7670 -2695 7685 -2670
rect 6000 -2710 6050 -2700
rect 7635 -2705 7685 -2695
rect 8175 -2670 8225 -2660
rect 8175 -2695 8190 -2670
rect 8210 -2695 8225 -2670
rect 8670 -2670 8685 -2640
rect 8730 -2670 8745 -2640
rect 8670 -2685 8745 -2670
rect 9305 -2640 9355 -2630
rect 9305 -2665 9320 -2640
rect 9340 -2665 9355 -2640
rect 9855 -2650 9870 -2625
rect 9890 -2650 9905 -2625
rect 10390 -2635 10405 -2605
rect 10450 -2635 10465 -2605
rect 11975 -2605 12050 -2590
rect 10390 -2650 10465 -2635
rect 10940 -2635 10990 -2625
rect 9855 -2660 9905 -2650
rect 10940 -2660 10955 -2635
rect 10975 -2660 10990 -2635
rect 9305 -2675 9355 -2665
rect 10940 -2670 10990 -2660
rect 11480 -2635 11530 -2625
rect 11480 -2660 11495 -2635
rect 11515 -2660 11530 -2635
rect 11975 -2635 11990 -2605
rect 12035 -2635 12050 -2605
rect 11975 -2650 12050 -2635
rect 12610 -2605 12660 -2595
rect 12610 -2630 12625 -2605
rect 12645 -2630 12660 -2605
rect 12610 -2640 12660 -2630
rect 11480 -2670 11530 -2660
rect 8175 -2705 8225 -2695
rect 4870 -2740 4920 -2730
rect 1565 -2775 1615 -2765
rect 130 -3890 180 -3880
rect 130 -3915 145 -3890
rect 165 -3915 180 -3890
rect 130 -3925 180 -3915
rect 3435 -3855 3485 -3845
rect 3435 -3880 3450 -3855
rect 3470 -3880 3485 -3855
rect 3435 -3890 3485 -3880
rect 1655 -4390 1705 -4380
rect 1655 -4415 1670 -4390
rect 1690 -4415 1705 -4390
rect 1655 -4425 1705 -4415
rect 6740 -3820 6790 -3810
rect 6740 -3845 6755 -3820
rect 6775 -3845 6790 -3820
rect 6740 -3855 6790 -3845
rect 4960 -4355 5010 -4345
rect 4960 -4380 4975 -4355
rect 4995 -4380 5010 -4355
rect 4960 -4390 5010 -4380
rect 10045 -3785 10095 -3775
rect 10045 -3810 10060 -3785
rect 10080 -3810 10095 -3785
rect 10045 -3820 10095 -3810
rect 2650 -4740 2700 -4730
rect 2650 -4765 2665 -4740
rect 2685 -4765 2700 -4740
rect 2650 -4775 2700 -4765
rect 8265 -4320 8315 -4310
rect 8265 -4345 8280 -4320
rect 8300 -4345 8315 -4320
rect 8265 -4355 8315 -4345
rect 13565 -4095 13615 -4085
rect 13135 -4135 13185 -4125
rect 13565 -4120 13580 -4095
rect 13600 -4120 13615 -4095
rect 13565 -4130 13615 -4120
rect 13135 -4160 13150 -4135
rect 13170 -4160 13185 -4135
rect 13135 -4170 13185 -4160
rect 5980 -4705 6030 -4695
rect 5980 -4730 5995 -4705
rect 6015 -4730 6030 -4705
rect 5980 -4740 6030 -4730
rect 11570 -4285 11620 -4275
rect 11570 -4310 11585 -4285
rect 11605 -4310 11620 -4285
rect 11570 -4320 11620 -4310
rect 9295 -4670 9345 -4660
rect 9295 -4695 9310 -4670
rect 9330 -4695 9345 -4670
rect 9295 -4705 9345 -4695
rect 80 -5150 130 -5140
rect 80 -5175 95 -5150
rect 115 -5175 130 -5150
rect 80 -5185 130 -5175
rect 3385 -5115 3435 -5105
rect 3385 -5140 3400 -5115
rect 3420 -5140 3435 -5115
rect 3385 -5150 3435 -5140
rect 6690 -5080 6740 -5070
rect 6690 -5105 6705 -5080
rect 6725 -5105 6740 -5080
rect 6690 -5115 6740 -5105
rect 9995 -5045 10045 -5035
rect 9995 -5070 10010 -5045
rect 10030 -5070 10045 -5045
rect 9995 -5080 10045 -5070
rect 9275 -6335 9325 -6325
rect 9275 -6360 9290 -6335
rect 9310 -6360 9325 -6335
rect 9275 -6370 9325 -6360
rect 6170 -6455 6220 -6445
rect 6170 -6480 6185 -6455
rect 6205 -6480 6220 -6455
rect 6170 -6490 6220 -6480
rect 2725 -6560 2775 -6550
rect 2725 -6585 2740 -6560
rect 2760 -6585 2775 -6560
rect 2725 -6595 2775 -6585
<< nsubdiff >>
rect 12595 -1655 12645 -1640
rect 9290 -1690 9340 -1675
rect 5985 -1725 6035 -1710
rect 2680 -1760 2730 -1745
rect 1550 -1790 1600 -1775
rect 1550 -1815 1565 -1790
rect 1585 -1815 1600 -1790
rect 2680 -1785 2695 -1760
rect 2715 -1785 2730 -1760
rect 2680 -1795 2730 -1785
rect 4855 -1755 4905 -1740
rect 4855 -1780 4870 -1755
rect 4890 -1780 4905 -1755
rect 5985 -1750 6000 -1725
rect 6020 -1750 6035 -1725
rect 5985 -1760 6035 -1750
rect 8160 -1720 8210 -1705
rect 8160 -1745 8175 -1720
rect 8195 -1745 8210 -1720
rect 9290 -1715 9305 -1690
rect 9325 -1715 9340 -1690
rect 9290 -1725 9340 -1715
rect 11465 -1685 11515 -1670
rect 11465 -1710 11480 -1685
rect 11500 -1710 11515 -1685
rect 12595 -1680 12610 -1655
rect 12630 -1680 12645 -1655
rect 12595 -1690 12645 -1680
rect 11465 -1720 11515 -1710
rect 8160 -1755 8210 -1745
rect 9815 -1755 9865 -1740
rect 4855 -1790 4905 -1780
rect 6510 -1790 6560 -1775
rect 9815 -1780 9830 -1755
rect 9850 -1780 9865 -1755
rect 1550 -1825 1600 -1815
rect 3205 -1825 3255 -1810
rect 6510 -1815 6525 -1790
rect 6545 -1815 6560 -1790
rect -100 -1860 -50 -1845
rect 3205 -1850 3220 -1825
rect 3240 -1850 3255 -1825
rect -100 -1885 -85 -1860
rect -65 -1885 -50 -1860
rect -100 -1895 -50 -1885
rect 490 -1875 540 -1860
rect 490 -1895 505 -1875
rect 525 -1895 540 -1875
rect 490 -1910 540 -1895
rect 985 -1870 1035 -1855
rect 3205 -1860 3255 -1850
rect 3795 -1840 3845 -1825
rect 3795 -1860 3810 -1840
rect 3830 -1860 3845 -1840
rect 985 -1895 1000 -1870
rect 1020 -1895 1035 -1870
rect 985 -1905 1035 -1895
rect 2075 -1875 2125 -1860
rect 3795 -1875 3845 -1860
rect 4290 -1835 4340 -1820
rect 6510 -1825 6560 -1815
rect 7100 -1805 7150 -1790
rect 7100 -1825 7115 -1805
rect 7135 -1825 7150 -1805
rect 4290 -1860 4305 -1835
rect 4325 -1860 4340 -1835
rect 4290 -1870 4340 -1860
rect 5380 -1840 5430 -1825
rect 7100 -1840 7150 -1825
rect 7595 -1800 7645 -1785
rect 9815 -1790 9865 -1780
rect 10405 -1770 10455 -1755
rect 10405 -1790 10420 -1770
rect 10440 -1790 10455 -1770
rect 7595 -1825 7610 -1800
rect 7630 -1825 7645 -1800
rect 7595 -1835 7645 -1825
rect 8685 -1805 8735 -1790
rect 10405 -1805 10455 -1790
rect 10900 -1765 10950 -1750
rect 10900 -1790 10915 -1765
rect 10935 -1790 10950 -1765
rect 10900 -1800 10950 -1790
rect 11990 -1770 12040 -1755
rect 11990 -1790 12005 -1770
rect 12025 -1790 12040 -1770
rect 11990 -1805 12040 -1790
rect 8685 -1825 8700 -1805
rect 8720 -1825 8735 -1805
rect 8685 -1840 8735 -1825
rect 5380 -1860 5395 -1840
rect 5415 -1860 5430 -1840
rect 5380 -1875 5430 -1860
rect 2075 -1895 2090 -1875
rect 2110 -1895 2125 -1875
rect 2075 -1910 2125 -1895
rect 10848 -2810 10898 -2795
rect 7543 -2845 7593 -2830
rect 4238 -2880 4288 -2865
rect 933 -2915 983 -2900
rect 115 -2940 165 -2925
rect 115 -2965 130 -2940
rect 150 -2965 165 -2940
rect 933 -2940 948 -2915
rect 968 -2940 983 -2915
rect 3420 -2905 3470 -2890
rect 3420 -2930 3435 -2905
rect 3455 -2930 3470 -2905
rect 4238 -2905 4253 -2880
rect 4273 -2905 4288 -2880
rect 6725 -2870 6775 -2855
rect 6725 -2895 6740 -2870
rect 6760 -2895 6775 -2870
rect 7543 -2870 7558 -2845
rect 7578 -2870 7593 -2845
rect 10030 -2835 10080 -2820
rect 10030 -2860 10045 -2835
rect 10065 -2860 10080 -2835
rect 10848 -2835 10863 -2810
rect 10883 -2835 10898 -2810
rect 10848 -2845 10898 -2835
rect 10030 -2870 10080 -2860
rect 7543 -2880 7593 -2870
rect 6725 -2905 6775 -2895
rect 4238 -2915 4288 -2905
rect 3420 -2940 3470 -2930
rect 933 -2950 983 -2940
rect 115 -2975 165 -2965
rect 2458 -3415 2508 -3400
rect 1640 -3440 1690 -3425
rect 1640 -3465 1655 -3440
rect 1675 -3465 1690 -3440
rect 2458 -3440 2473 -3415
rect 2493 -3440 2508 -3415
rect 2458 -3450 2508 -3440
rect 1640 -3475 1690 -3465
rect 928 -3510 978 -3495
rect 928 -3535 943 -3510
rect 963 -3535 978 -3510
rect 928 -3545 978 -3535
rect 5763 -3380 5813 -3365
rect 4945 -3405 4995 -3390
rect 4945 -3430 4960 -3405
rect 4980 -3430 4995 -3405
rect 5763 -3405 5778 -3380
rect 5798 -3405 5813 -3380
rect 5763 -3415 5813 -3405
rect 4945 -3440 4995 -3430
rect 4233 -3475 4283 -3460
rect 4233 -3500 4248 -3475
rect 4268 -3500 4283 -3475
rect 4233 -3510 4283 -3500
rect 9068 -3345 9118 -3330
rect 8250 -3370 8300 -3355
rect 8250 -3395 8265 -3370
rect 8285 -3395 8300 -3370
rect 9068 -3370 9083 -3345
rect 9103 -3370 9118 -3345
rect 9068 -3380 9118 -3370
rect 8250 -3405 8300 -3395
rect 7538 -3440 7588 -3425
rect 7538 -3465 7553 -3440
rect 7573 -3465 7588 -3440
rect 7538 -3475 7588 -3465
rect 2720 -3710 2770 -3695
rect 2720 -3735 2735 -3710
rect 2755 -3735 2770 -3710
rect 2720 -3745 2770 -3735
rect 2453 -4010 2503 -3995
rect 2453 -4035 2468 -4010
rect 2488 -4035 2503 -4010
rect 2453 -4045 2503 -4035
rect 883 -4175 933 -4160
rect 65 -4200 115 -4185
rect 65 -4225 80 -4200
rect 100 -4225 115 -4200
rect 883 -4200 898 -4175
rect 918 -4200 933 -4175
rect 883 -4210 933 -4200
rect 65 -4235 115 -4225
rect 13635 -3065 13685 -3050
rect 13635 -3090 13650 -3065
rect 13670 -3090 13685 -3065
rect 13205 -3105 13255 -3090
rect 13635 -3100 13685 -3090
rect 13205 -3130 13220 -3105
rect 13240 -3130 13255 -3105
rect 13205 -3140 13255 -3130
rect 12373 -3310 12423 -3295
rect 11555 -3335 11605 -3320
rect 11555 -3360 11570 -3335
rect 11590 -3360 11605 -3335
rect 12373 -3335 12388 -3310
rect 12408 -3335 12423 -3310
rect 12373 -3345 12423 -3335
rect 11555 -3370 11605 -3360
rect 10843 -3405 10893 -3390
rect 10843 -3430 10858 -3405
rect 10878 -3430 10893 -3405
rect 10843 -3440 10893 -3430
rect 6050 -3675 6100 -3660
rect 6050 -3700 6065 -3675
rect 6085 -3700 6100 -3675
rect 6050 -3710 6100 -3700
rect 5758 -3975 5808 -3960
rect 5758 -4000 5773 -3975
rect 5793 -4000 5808 -3975
rect 5758 -4010 5808 -4000
rect 4188 -4140 4238 -4125
rect 3370 -4165 3420 -4150
rect 3370 -4190 3385 -4165
rect 3405 -4190 3420 -4165
rect 4188 -4165 4203 -4140
rect 4223 -4165 4238 -4140
rect 4188 -4175 4238 -4165
rect 3370 -4200 3420 -4190
rect 9365 -3640 9415 -3625
rect 9365 -3665 9380 -3640
rect 9400 -3665 9415 -3640
rect 9365 -3675 9415 -3665
rect 9063 -3940 9113 -3925
rect 9063 -3965 9078 -3940
rect 9098 -3965 9113 -3940
rect 9063 -3975 9113 -3965
rect 7493 -4105 7543 -4090
rect 6675 -4130 6725 -4115
rect 6675 -4155 6690 -4130
rect 6710 -4155 6725 -4130
rect 7493 -4130 7508 -4105
rect 7528 -4130 7543 -4105
rect 7493 -4140 7543 -4130
rect 6675 -4165 6725 -4155
rect 878 -4770 928 -4755
rect 878 -4795 893 -4770
rect 913 -4795 928 -4770
rect 12368 -3905 12418 -3890
rect 12368 -3930 12383 -3905
rect 12403 -3930 12418 -3905
rect 12368 -3940 12418 -3930
rect 10798 -4070 10848 -4055
rect 9980 -4095 10030 -4080
rect 9980 -4120 9995 -4095
rect 10015 -4120 10030 -4095
rect 10798 -4095 10813 -4070
rect 10833 -4095 10848 -4070
rect 10798 -4105 10848 -4095
rect 9980 -4130 10030 -4120
rect 4183 -4735 4233 -4720
rect 4183 -4760 4198 -4735
rect 4218 -4760 4233 -4735
rect 7488 -4700 7538 -4685
rect 7488 -4725 7503 -4700
rect 7523 -4725 7538 -4700
rect 10793 -4665 10843 -4650
rect 10793 -4690 10808 -4665
rect 10828 -4690 10843 -4665
rect 10793 -4700 10843 -4690
rect 7488 -4735 7538 -4725
rect 4183 -4770 4233 -4760
rect 878 -4805 928 -4795
rect 9345 -5305 9395 -5290
rect 9345 -5330 9360 -5305
rect 9380 -5330 9395 -5305
rect 9345 -5340 9395 -5330
rect 6240 -5425 6290 -5410
rect 6240 -5450 6255 -5425
rect 6275 -5450 6290 -5425
rect 6240 -5460 6290 -5450
rect 2795 -5530 2845 -5515
rect 2795 -5555 2810 -5530
rect 2830 -5555 2845 -5530
rect 2795 -5565 2845 -5555
<< psubdiffcont >>
rect -45 -2755 -25 -2730
rect 490 -2740 535 -2710
rect 1040 -2765 1060 -2740
rect 1580 -2765 1600 -2740
rect 2075 -2740 2120 -2710
rect 2710 -2735 2730 -2710
rect 3260 -2720 3280 -2695
rect 3795 -2705 3840 -2675
rect 4345 -2730 4365 -2705
rect 4885 -2730 4905 -2705
rect 5380 -2705 5425 -2675
rect 6015 -2700 6035 -2675
rect 6565 -2685 6585 -2660
rect 7100 -2670 7145 -2640
rect 7650 -2695 7670 -2670
rect 8190 -2695 8210 -2670
rect 8685 -2670 8730 -2640
rect 9320 -2665 9340 -2640
rect 9870 -2650 9890 -2625
rect 10405 -2635 10450 -2605
rect 10955 -2660 10975 -2635
rect 11495 -2660 11515 -2635
rect 11990 -2635 12035 -2605
rect 12625 -2630 12645 -2605
rect 145 -3915 165 -3890
rect 3450 -3880 3470 -3855
rect 1670 -4415 1690 -4390
rect 6755 -3845 6775 -3820
rect 4975 -4380 4995 -4355
rect 10060 -3810 10080 -3785
rect 2665 -4765 2685 -4740
rect 8280 -4345 8300 -4320
rect 13580 -4120 13600 -4095
rect 13150 -4160 13170 -4135
rect 5995 -4730 6015 -4705
rect 11585 -4310 11605 -4285
rect 9310 -4695 9330 -4670
rect 95 -5175 115 -5150
rect 3400 -5140 3420 -5115
rect 6705 -5105 6725 -5080
rect 10010 -5070 10030 -5045
rect 9290 -6360 9310 -6335
rect 6185 -6480 6205 -6455
rect 2740 -6585 2760 -6560
<< nsubdiffcont >>
rect 1565 -1815 1585 -1790
rect 2695 -1785 2715 -1760
rect 4870 -1780 4890 -1755
rect 6000 -1750 6020 -1725
rect 8175 -1745 8195 -1720
rect 9305 -1715 9325 -1690
rect 11480 -1710 11500 -1685
rect 12610 -1680 12630 -1655
rect 9830 -1780 9850 -1755
rect 6525 -1815 6545 -1790
rect 3220 -1850 3240 -1825
rect -85 -1885 -65 -1860
rect 505 -1895 525 -1875
rect 3810 -1860 3830 -1840
rect 1000 -1895 1020 -1870
rect 7115 -1825 7135 -1805
rect 4305 -1860 4325 -1835
rect 10420 -1790 10440 -1770
rect 7610 -1825 7630 -1800
rect 10915 -1790 10935 -1765
rect 12005 -1790 12025 -1770
rect 8700 -1825 8720 -1805
rect 5395 -1860 5415 -1840
rect 2090 -1895 2110 -1875
rect 130 -2965 150 -2940
rect 948 -2940 968 -2915
rect 3435 -2930 3455 -2905
rect 4253 -2905 4273 -2880
rect 6740 -2895 6760 -2870
rect 7558 -2870 7578 -2845
rect 10045 -2860 10065 -2835
rect 10863 -2835 10883 -2810
rect 1655 -3465 1675 -3440
rect 2473 -3440 2493 -3415
rect 943 -3535 963 -3510
rect 4960 -3430 4980 -3405
rect 5778 -3405 5798 -3380
rect 4248 -3500 4268 -3475
rect 8265 -3395 8285 -3370
rect 9083 -3370 9103 -3345
rect 7553 -3465 7573 -3440
rect 2735 -3735 2755 -3710
rect 2468 -4035 2488 -4010
rect 80 -4225 100 -4200
rect 898 -4200 918 -4175
rect 13650 -3090 13670 -3065
rect 13220 -3130 13240 -3105
rect 11570 -3360 11590 -3335
rect 12388 -3335 12408 -3310
rect 10858 -3430 10878 -3405
rect 6065 -3700 6085 -3675
rect 5773 -4000 5793 -3975
rect 3385 -4190 3405 -4165
rect 4203 -4165 4223 -4140
rect 9380 -3665 9400 -3640
rect 9078 -3965 9098 -3940
rect 6690 -4155 6710 -4130
rect 7508 -4130 7528 -4105
rect 893 -4795 913 -4770
rect 12383 -3930 12403 -3905
rect 9995 -4120 10015 -4095
rect 10813 -4095 10833 -4070
rect 4198 -4760 4218 -4735
rect 7503 -4725 7523 -4700
rect 10808 -4690 10828 -4665
rect 9360 -5330 9380 -5305
rect 6255 -5450 6275 -5425
rect 2810 -5555 2830 -5530
<< poly >>
rect 165 -1965 180 -1930
rect 250 -1965 265 -1930
rect 660 -1950 675 -1910
rect 750 -1950 765 -1910
rect 165 -2210 180 -2165
rect 120 -2220 180 -2210
rect 120 -2245 130 -2220
rect 160 -2245 180 -2220
rect 120 -2255 180 -2245
rect 165 -2465 180 -2255
rect 250 -2370 265 -2165
rect 1255 -1975 1270 -1940
rect 1335 -1975 1350 -1940
rect 1800 -1975 1815 -1935
rect 2245 -1950 2260 -1910
rect 2335 -1950 2350 -1910
rect 2930 -1945 2945 -1905
rect 3470 -1930 3485 -1895
rect 3555 -1930 3570 -1895
rect 3965 -1915 3980 -1875
rect 4055 -1915 4070 -1875
rect 1255 -2220 1270 -2175
rect 1205 -2230 1270 -2220
rect 1205 -2255 1215 -2230
rect 1245 -2255 1270 -2230
rect 1205 -2265 1270 -2255
rect 210 -2380 265 -2370
rect 210 -2405 220 -2380
rect 240 -2405 265 -2380
rect 660 -2385 675 -2350
rect 210 -2415 265 -2405
rect 620 -2390 675 -2385
rect 620 -2410 630 -2390
rect 650 -2410 675 -2390
rect 620 -2415 675 -2410
rect 250 -2465 265 -2415
rect 660 -2575 675 -2415
rect 750 -2465 765 -2350
rect 710 -2470 765 -2465
rect 710 -2490 720 -2470
rect 740 -2490 765 -2470
rect 1255 -2475 1270 -2265
rect 1335 -2380 1350 -2175
rect 1800 -2355 1815 -2175
rect 2930 -2325 2945 -2145
rect 3470 -2175 3485 -2130
rect 3425 -2185 3485 -2175
rect 3425 -2210 3435 -2185
rect 3465 -2210 3485 -2185
rect 3425 -2220 3485 -2210
rect 2855 -2340 2945 -2325
rect 1295 -2390 1350 -2380
rect 1295 -2415 1305 -2390
rect 1325 -2415 1350 -2390
rect 1725 -2370 1815 -2355
rect 1725 -2395 1750 -2370
rect 1780 -2395 1815 -2370
rect 2245 -2385 2260 -2350
rect 1725 -2405 1815 -2395
rect 1295 -2425 1350 -2415
rect 1335 -2475 1350 -2425
rect 710 -2495 765 -2490
rect 750 -2575 765 -2495
rect 165 -2685 180 -2665
rect 250 -2685 265 -2665
rect 1800 -2575 1815 -2405
rect 2205 -2390 2260 -2385
rect 2205 -2410 2215 -2390
rect 2235 -2410 2260 -2390
rect 2205 -2415 2260 -2410
rect 2245 -2575 2260 -2415
rect 2335 -2465 2350 -2350
rect 2855 -2365 2880 -2340
rect 2910 -2365 2945 -2340
rect 2855 -2375 2945 -2365
rect 2295 -2470 2350 -2465
rect 2295 -2490 2305 -2470
rect 2325 -2490 2350 -2470
rect 2295 -2495 2350 -2490
rect 2335 -2575 2350 -2495
rect 2930 -2545 2945 -2375
rect 3470 -2430 3485 -2220
rect 3555 -2335 3570 -2130
rect 4560 -1940 4575 -1905
rect 4640 -1940 4655 -1905
rect 5105 -1940 5120 -1900
rect 5550 -1915 5565 -1875
rect 5640 -1915 5655 -1875
rect 6235 -1910 6250 -1870
rect 6775 -1895 6790 -1860
rect 6860 -1895 6875 -1860
rect 7270 -1880 7285 -1840
rect 7360 -1880 7375 -1840
rect 4560 -2185 4575 -2140
rect 4510 -2195 4575 -2185
rect 4510 -2220 4520 -2195
rect 4550 -2220 4575 -2195
rect 4510 -2230 4575 -2220
rect 3515 -2345 3570 -2335
rect 3515 -2370 3525 -2345
rect 3545 -2370 3570 -2345
rect 3965 -2350 3980 -2315
rect 3515 -2380 3570 -2370
rect 3925 -2355 3980 -2350
rect 3925 -2375 3935 -2355
rect 3955 -2375 3980 -2355
rect 3925 -2380 3980 -2375
rect 3555 -2430 3570 -2380
rect 3965 -2540 3980 -2380
rect 4055 -2430 4070 -2315
rect 4015 -2435 4070 -2430
rect 4015 -2455 4025 -2435
rect 4045 -2455 4070 -2435
rect 4560 -2440 4575 -2230
rect 4640 -2345 4655 -2140
rect 5105 -2320 5120 -2140
rect 6235 -2290 6250 -2110
rect 6775 -2140 6790 -2095
rect 6730 -2150 6790 -2140
rect 6730 -2175 6740 -2150
rect 6770 -2175 6790 -2150
rect 6730 -2185 6790 -2175
rect 6160 -2305 6250 -2290
rect 4600 -2355 4655 -2345
rect 4600 -2380 4610 -2355
rect 4630 -2380 4655 -2355
rect 5030 -2335 5120 -2320
rect 5030 -2360 5055 -2335
rect 5085 -2360 5120 -2335
rect 5550 -2350 5565 -2315
rect 5030 -2370 5120 -2360
rect 4600 -2390 4655 -2380
rect 4640 -2440 4655 -2390
rect 4015 -2460 4070 -2455
rect 4055 -2540 4070 -2460
rect 2930 -2660 2945 -2645
rect 3470 -2650 3485 -2630
rect 3555 -2650 3570 -2630
rect 5105 -2540 5120 -2370
rect 5510 -2355 5565 -2350
rect 5510 -2375 5520 -2355
rect 5540 -2375 5565 -2355
rect 5510 -2380 5565 -2375
rect 5550 -2540 5565 -2380
rect 5640 -2430 5655 -2315
rect 6160 -2330 6185 -2305
rect 6215 -2330 6250 -2305
rect 6160 -2340 6250 -2330
rect 5600 -2435 5655 -2430
rect 5600 -2455 5610 -2435
rect 5630 -2455 5655 -2435
rect 5600 -2460 5655 -2455
rect 5640 -2540 5655 -2460
rect 6235 -2510 6250 -2340
rect 6775 -2395 6790 -2185
rect 6860 -2300 6875 -2095
rect 7865 -1905 7880 -1870
rect 7945 -1905 7960 -1870
rect 8410 -1905 8425 -1865
rect 8855 -1880 8870 -1840
rect 8945 -1880 8960 -1840
rect 9540 -1875 9555 -1835
rect 10080 -1860 10095 -1825
rect 10165 -1860 10180 -1825
rect 10575 -1845 10590 -1805
rect 10665 -1845 10680 -1805
rect 7865 -2150 7880 -2105
rect 7815 -2160 7880 -2150
rect 7815 -2185 7825 -2160
rect 7855 -2185 7880 -2160
rect 7815 -2195 7880 -2185
rect 6820 -2310 6875 -2300
rect 6820 -2335 6830 -2310
rect 6850 -2335 6875 -2310
rect 7270 -2315 7285 -2280
rect 6820 -2345 6875 -2335
rect 7230 -2320 7285 -2315
rect 7230 -2340 7240 -2320
rect 7260 -2340 7285 -2320
rect 7230 -2345 7285 -2340
rect 6860 -2395 6875 -2345
rect 7270 -2505 7285 -2345
rect 7360 -2395 7375 -2280
rect 7320 -2400 7375 -2395
rect 7320 -2420 7330 -2400
rect 7350 -2420 7375 -2400
rect 7865 -2405 7880 -2195
rect 7945 -2310 7960 -2105
rect 8410 -2285 8425 -2105
rect 9540 -2255 9555 -2075
rect 10080 -2105 10095 -2060
rect 10035 -2115 10095 -2105
rect 10035 -2140 10045 -2115
rect 10075 -2140 10095 -2115
rect 10035 -2150 10095 -2140
rect 9465 -2270 9555 -2255
rect 7905 -2320 7960 -2310
rect 7905 -2345 7915 -2320
rect 7935 -2345 7960 -2320
rect 8335 -2300 8425 -2285
rect 8335 -2325 8360 -2300
rect 8390 -2325 8425 -2300
rect 8855 -2315 8870 -2280
rect 8335 -2335 8425 -2325
rect 7905 -2355 7960 -2345
rect 7945 -2405 7960 -2355
rect 7320 -2425 7375 -2420
rect 7360 -2505 7375 -2425
rect 6235 -2625 6250 -2610
rect 6775 -2615 6790 -2595
rect 6860 -2615 6875 -2595
rect 8410 -2505 8425 -2335
rect 8815 -2320 8870 -2315
rect 8815 -2340 8825 -2320
rect 8845 -2340 8870 -2320
rect 8815 -2345 8870 -2340
rect 8855 -2505 8870 -2345
rect 8945 -2395 8960 -2280
rect 9465 -2295 9490 -2270
rect 9520 -2295 9555 -2270
rect 9465 -2305 9555 -2295
rect 8905 -2400 8960 -2395
rect 8905 -2420 8915 -2400
rect 8935 -2420 8960 -2400
rect 8905 -2425 8960 -2420
rect 8945 -2505 8960 -2425
rect 9540 -2475 9555 -2305
rect 10080 -2360 10095 -2150
rect 10165 -2265 10180 -2060
rect 11170 -1870 11185 -1835
rect 11250 -1870 11265 -1835
rect 11715 -1870 11730 -1830
rect 12160 -1845 12175 -1805
rect 12250 -1845 12265 -1805
rect 12845 -1840 12860 -1800
rect 11170 -2115 11185 -2070
rect 11120 -2125 11185 -2115
rect 11120 -2150 11130 -2125
rect 11160 -2150 11185 -2125
rect 11120 -2160 11185 -2150
rect 10125 -2275 10180 -2265
rect 10125 -2300 10135 -2275
rect 10155 -2300 10180 -2275
rect 10575 -2280 10590 -2245
rect 10125 -2310 10180 -2300
rect 10535 -2285 10590 -2280
rect 10535 -2305 10545 -2285
rect 10565 -2305 10590 -2285
rect 10535 -2310 10590 -2305
rect 10165 -2360 10180 -2310
rect 10575 -2470 10590 -2310
rect 10665 -2360 10680 -2245
rect 10625 -2365 10680 -2360
rect 10625 -2385 10635 -2365
rect 10655 -2385 10680 -2365
rect 11170 -2370 11185 -2160
rect 11250 -2275 11265 -2070
rect 11715 -2250 11730 -2070
rect 12845 -2220 12860 -2040
rect 12770 -2235 12860 -2220
rect 11210 -2285 11265 -2275
rect 11210 -2310 11220 -2285
rect 11240 -2310 11265 -2285
rect 11640 -2265 11730 -2250
rect 11640 -2290 11665 -2265
rect 11695 -2290 11730 -2265
rect 12160 -2280 12175 -2245
rect 11640 -2300 11730 -2290
rect 11210 -2320 11265 -2310
rect 11250 -2370 11265 -2320
rect 10625 -2390 10680 -2385
rect 10665 -2470 10680 -2390
rect 9540 -2590 9555 -2575
rect 10080 -2580 10095 -2560
rect 10165 -2580 10180 -2560
rect 11715 -2470 11730 -2300
rect 12120 -2285 12175 -2280
rect 12120 -2305 12130 -2285
rect 12150 -2305 12175 -2285
rect 12120 -2310 12175 -2305
rect 12160 -2470 12175 -2310
rect 12250 -2360 12265 -2245
rect 12770 -2260 12795 -2235
rect 12825 -2260 12860 -2235
rect 12770 -2270 12860 -2260
rect 12210 -2365 12265 -2360
rect 12210 -2385 12220 -2365
rect 12240 -2385 12265 -2365
rect 12210 -2390 12265 -2385
rect 12250 -2470 12265 -2390
rect 12845 -2440 12860 -2270
rect 12845 -2555 12860 -2540
rect 10575 -2590 10590 -2570
rect 10665 -2590 10680 -2570
rect 11170 -2590 11185 -2570
rect 11250 -2590 11265 -2570
rect 11715 -2585 11730 -2570
rect 12160 -2590 12175 -2570
rect 12250 -2590 12265 -2570
rect 7270 -2625 7285 -2605
rect 7360 -2625 7375 -2605
rect 7865 -2625 7880 -2605
rect 7945 -2625 7960 -2605
rect 8410 -2620 8425 -2605
rect 8855 -2625 8870 -2605
rect 8945 -2625 8960 -2605
rect 3965 -2660 3980 -2640
rect 4055 -2660 4070 -2640
rect 4560 -2660 4575 -2640
rect 4640 -2660 4655 -2640
rect 5105 -2655 5120 -2640
rect 5550 -2660 5565 -2640
rect 5640 -2660 5655 -2640
rect 660 -2695 675 -2675
rect 750 -2695 765 -2675
rect 1255 -2695 1270 -2675
rect 1335 -2695 1350 -2675
rect 1800 -2690 1815 -2675
rect 2245 -2695 2260 -2675
rect 2335 -2695 2350 -2675
rect 10895 -2885 10910 -2870
rect 7590 -2920 7605 -2905
rect 4285 -2955 4300 -2940
rect 980 -2990 995 -2975
rect 365 -3095 730 -3080
rect 3670 -3060 4035 -3045
rect 6975 -3025 7340 -3010
rect 10280 -2990 10645 -2975
rect 10280 -3020 10295 -2990
rect 10620 -2995 10645 -2990
rect 10895 -2995 10910 -2985
rect 10620 -3010 10910 -2995
rect 6975 -3055 6990 -3025
rect 7315 -3030 7340 -3025
rect 7590 -3030 7605 -3020
rect 7315 -3045 7605 -3030
rect 3670 -3090 3685 -3060
rect 4010 -3065 4035 -3060
rect 4285 -3065 4300 -3055
rect 4010 -3080 4300 -3065
rect 365 -3125 380 -3095
rect 705 -3100 730 -3095
rect 980 -3100 995 -3090
rect 705 -3115 995 -3100
rect 685 -3180 995 -3160
rect 365 -3505 380 -3325
rect 290 -3520 380 -3505
rect 290 -3545 315 -3520
rect 345 -3545 380 -3520
rect 290 -3555 380 -3545
rect 685 -3555 710 -3180
rect 980 -3190 995 -3180
rect 3990 -3145 4300 -3125
rect 980 -3310 995 -3290
rect 2505 -3490 2520 -3460
rect 3670 -3470 3685 -3290
rect 3595 -3485 3685 -3470
rect 365 -3725 380 -3555
rect 675 -3560 715 -3555
rect 675 -3585 685 -3560
rect 705 -3585 715 -3560
rect 975 -3585 990 -3565
rect 675 -3590 715 -3585
rect 685 -3710 710 -3590
rect 1890 -3595 2285 -3580
rect 3595 -3510 3620 -3485
rect 3650 -3510 3685 -3485
rect 3595 -3520 3685 -3510
rect 3990 -3520 4015 -3145
rect 4285 -3155 4300 -3145
rect 7295 -3110 7605 -3090
rect 4285 -3275 4300 -3255
rect 5810 -3455 5825 -3425
rect 6975 -3435 6990 -3255
rect 6900 -3450 6990 -3435
rect 1890 -3625 1905 -3595
rect 2255 -3600 2285 -3595
rect 2505 -3600 2520 -3590
rect 2255 -3615 2520 -3600
rect 975 -3710 990 -3685
rect 685 -3730 990 -3710
rect 975 -3785 990 -3770
rect 365 -3835 380 -3825
rect 365 -3850 790 -3835
rect 775 -3910 790 -3850
rect 2210 -3680 2520 -3660
rect 975 -3910 990 -3885
rect 775 -3925 990 -3910
rect 1890 -4005 1905 -3825
rect 1815 -4020 1905 -4005
rect 1815 -4045 1840 -4020
rect 1870 -4045 1905 -4020
rect 1815 -4055 1905 -4045
rect 2210 -4055 2235 -3680
rect 2505 -3690 2520 -3680
rect 3670 -3690 3685 -3520
rect 3980 -3525 4020 -3520
rect 3980 -3550 3990 -3525
rect 4010 -3550 4020 -3525
rect 4280 -3550 4295 -3530
rect 3980 -3555 4020 -3550
rect 3990 -3675 4015 -3555
rect 5195 -3560 5590 -3545
rect 6900 -3475 6925 -3450
rect 6955 -3475 6990 -3450
rect 6900 -3485 6990 -3475
rect 7295 -3485 7320 -3110
rect 7590 -3120 7605 -3110
rect 10600 -3075 10910 -3055
rect 7590 -3240 7605 -3220
rect 9115 -3420 9130 -3390
rect 10280 -3400 10295 -3220
rect 10205 -3415 10295 -3400
rect 5195 -3590 5210 -3560
rect 5560 -3565 5590 -3560
rect 5810 -3565 5825 -3555
rect 5560 -3580 5825 -3565
rect 4280 -3675 4295 -3650
rect 3990 -3695 4295 -3675
rect 4280 -3750 4295 -3735
rect 2505 -3810 2520 -3790
rect 3670 -3800 3685 -3790
rect 3670 -3815 4095 -3800
rect 4080 -3875 4095 -3815
rect 5515 -3645 5825 -3625
rect 4280 -3875 4295 -3850
rect 4080 -3890 4295 -3875
rect 2900 -3915 2915 -3890
rect 930 -4250 945 -4220
rect 1890 -4225 1905 -4055
rect 2200 -4060 2240 -4055
rect 2200 -4085 2210 -4060
rect 2230 -4085 2240 -4060
rect 2500 -4085 2515 -4065
rect 2200 -4090 2240 -4085
rect 2210 -4210 2235 -4090
rect 2500 -4210 2515 -4185
rect 315 -4355 825 -4340
rect 2210 -4230 2515 -4210
rect 2500 -4285 2515 -4270
rect 1890 -4335 1905 -4325
rect 1890 -4350 2315 -4335
rect 315 -4385 330 -4355
rect 800 -4360 825 -4355
rect 930 -4360 945 -4350
rect 800 -4375 945 -4360
rect 635 -4440 945 -4420
rect 2300 -4410 2315 -4350
rect 5195 -3970 5210 -3790
rect 5120 -3985 5210 -3970
rect 5120 -4010 5145 -3985
rect 5175 -4010 5210 -3985
rect 5120 -4020 5210 -4010
rect 5515 -4020 5540 -3645
rect 5810 -3655 5825 -3645
rect 6975 -3655 6990 -3485
rect 7285 -3490 7325 -3485
rect 7285 -3515 7295 -3490
rect 7315 -3515 7325 -3490
rect 7585 -3515 7600 -3495
rect 7285 -3520 7325 -3515
rect 7295 -3640 7320 -3520
rect 8500 -3525 8895 -3510
rect 10205 -3440 10230 -3415
rect 10260 -3440 10295 -3415
rect 10205 -3450 10295 -3440
rect 10600 -3450 10625 -3075
rect 10895 -3085 10910 -3075
rect 10895 -3205 10910 -3185
rect 13815 -3270 13830 -3245
rect 13385 -3310 13400 -3285
rect 12420 -3385 12435 -3355
rect 8500 -3555 8515 -3525
rect 8865 -3530 8895 -3525
rect 9115 -3530 9130 -3520
rect 8865 -3545 9130 -3530
rect 7585 -3640 7600 -3615
rect 7295 -3660 7600 -3640
rect 7585 -3715 7600 -3700
rect 5810 -3775 5825 -3755
rect 6975 -3765 6990 -3755
rect 6975 -3780 7400 -3765
rect 7385 -3840 7400 -3780
rect 8820 -3610 9130 -3590
rect 7585 -3840 7600 -3815
rect 7385 -3855 7600 -3840
rect 6230 -3880 6245 -3855
rect 4235 -4215 4250 -4185
rect 5195 -4190 5210 -4020
rect 5505 -4025 5545 -4020
rect 5505 -4050 5515 -4025
rect 5535 -4050 5545 -4025
rect 5805 -4050 5820 -4030
rect 5505 -4055 5545 -4050
rect 5515 -4175 5540 -4055
rect 5805 -4175 5820 -4150
rect 2900 -4385 2915 -4315
rect 3620 -4320 4130 -4305
rect 5515 -4195 5820 -4175
rect 5805 -4250 5820 -4235
rect 5195 -4300 5210 -4290
rect 5195 -4315 5620 -4300
rect 3620 -4350 3635 -4320
rect 4105 -4325 4130 -4320
rect 4235 -4325 4250 -4315
rect 4105 -4340 4250 -4325
rect 2500 -4410 2515 -4385
rect 2300 -4425 2515 -4410
rect 2860 -4395 2915 -4385
rect 2860 -4415 2870 -4395
rect 2890 -4415 2915 -4395
rect 2860 -4425 2915 -4415
rect 315 -4765 330 -4585
rect 240 -4780 330 -4765
rect 240 -4805 265 -4780
rect 295 -4805 330 -4780
rect 240 -4815 330 -4805
rect 635 -4815 660 -4440
rect 930 -4450 945 -4440
rect 2900 -4515 2915 -4425
rect 930 -4570 945 -4550
rect 3940 -4405 4250 -4385
rect 5605 -4375 5620 -4315
rect 8500 -3935 8515 -3755
rect 8425 -3950 8515 -3935
rect 8425 -3975 8450 -3950
rect 8480 -3975 8515 -3950
rect 8425 -3985 8515 -3975
rect 8820 -3985 8845 -3610
rect 9115 -3620 9130 -3610
rect 10280 -3620 10295 -3450
rect 10590 -3455 10630 -3450
rect 10590 -3480 10600 -3455
rect 10620 -3480 10630 -3455
rect 10890 -3480 10905 -3460
rect 10590 -3485 10630 -3480
rect 10600 -3605 10625 -3485
rect 11805 -3490 12200 -3475
rect 11805 -3520 11820 -3490
rect 12170 -3495 12200 -3490
rect 12420 -3495 12435 -3485
rect 12170 -3510 12435 -3495
rect 10890 -3605 10905 -3580
rect 10600 -3625 10905 -3605
rect 10890 -3680 10905 -3665
rect 9115 -3740 9130 -3720
rect 10280 -3730 10295 -3720
rect 10280 -3745 10705 -3730
rect 10690 -3805 10705 -3745
rect 12125 -3575 12435 -3555
rect 10890 -3805 10905 -3780
rect 10690 -3820 10905 -3805
rect 9545 -3845 9560 -3820
rect 7540 -4180 7555 -4150
rect 8500 -4155 8515 -3985
rect 8810 -3990 8850 -3985
rect 8810 -4015 8820 -3990
rect 8840 -4015 8850 -3990
rect 9110 -4015 9125 -3995
rect 8810 -4020 8850 -4015
rect 8820 -4140 8845 -4020
rect 9110 -4140 9125 -4115
rect 6230 -4350 6245 -4280
rect 6925 -4285 7435 -4270
rect 8820 -4160 9125 -4140
rect 9110 -4215 9125 -4200
rect 8500 -4265 8515 -4255
rect 8500 -4280 8925 -4265
rect 6925 -4315 6940 -4285
rect 7410 -4290 7435 -4285
rect 7540 -4290 7555 -4280
rect 7410 -4305 7555 -4290
rect 5805 -4375 5820 -4350
rect 5605 -4390 5820 -4375
rect 6190 -4360 6245 -4350
rect 6190 -4380 6200 -4360
rect 6220 -4380 6245 -4360
rect 6190 -4390 6245 -4380
rect 2900 -4740 2915 -4715
rect 3620 -4730 3635 -4550
rect 3545 -4745 3635 -4730
rect 3545 -4770 3570 -4745
rect 3600 -4770 3635 -4745
rect 3545 -4780 3635 -4770
rect 3940 -4780 3965 -4405
rect 4235 -4415 4250 -4405
rect 6230 -4480 6245 -4390
rect 4235 -4535 4250 -4515
rect 7245 -4370 7555 -4350
rect 8910 -4340 8925 -4280
rect 11805 -3900 11820 -3720
rect 11730 -3915 11820 -3900
rect 11730 -3940 11755 -3915
rect 11785 -3940 11820 -3915
rect 11730 -3950 11820 -3940
rect 12125 -3950 12150 -3575
rect 12420 -3585 12435 -3575
rect 12420 -3705 12435 -3685
rect 13385 -3780 13400 -3710
rect 13815 -3740 13830 -3670
rect 13775 -3750 13830 -3740
rect 13775 -3770 13785 -3750
rect 13805 -3770 13830 -3750
rect 13775 -3780 13830 -3770
rect 13345 -3790 13400 -3780
rect 13345 -3810 13355 -3790
rect 13375 -3810 13400 -3790
rect 13345 -3820 13400 -3810
rect 13385 -3910 13400 -3820
rect 13815 -3870 13830 -3780
rect 10845 -4145 10860 -4115
rect 11805 -4120 11820 -3950
rect 12115 -3955 12155 -3950
rect 12115 -3980 12125 -3955
rect 12145 -3980 12155 -3955
rect 12415 -3980 12430 -3960
rect 12115 -3985 12155 -3980
rect 12125 -4105 12150 -3985
rect 12415 -4105 12430 -4080
rect 9545 -4315 9560 -4245
rect 10230 -4250 10740 -4235
rect 12125 -4125 12430 -4105
rect 13815 -4095 13830 -4070
rect 13385 -4135 13400 -4110
rect 12415 -4180 12430 -4165
rect 11805 -4230 11820 -4220
rect 11805 -4245 12230 -4230
rect 10230 -4280 10245 -4250
rect 10715 -4255 10740 -4250
rect 10845 -4255 10860 -4245
rect 10715 -4270 10860 -4255
rect 9110 -4340 9125 -4315
rect 8910 -4355 9125 -4340
rect 9505 -4325 9560 -4315
rect 9505 -4345 9515 -4325
rect 9535 -4345 9560 -4325
rect 9505 -4355 9560 -4345
rect 6230 -4705 6245 -4680
rect 6925 -4695 6940 -4515
rect 6850 -4710 6940 -4695
rect 6850 -4735 6875 -4710
rect 6905 -4735 6940 -4710
rect 6850 -4745 6940 -4735
rect 7245 -4745 7270 -4370
rect 7540 -4380 7555 -4370
rect 9545 -4445 9560 -4355
rect 7540 -4500 7555 -4480
rect 10550 -4335 10860 -4315
rect 12215 -4305 12230 -4245
rect 12415 -4305 12430 -4280
rect 12215 -4320 12430 -4305
rect 9545 -4670 9560 -4645
rect 10230 -4660 10245 -4480
rect 10155 -4675 10245 -4660
rect 10155 -4700 10180 -4675
rect 10210 -4700 10245 -4675
rect 10155 -4710 10245 -4700
rect 10550 -4710 10575 -4335
rect 10845 -4345 10860 -4335
rect 10845 -4465 10860 -4445
rect 315 -4985 330 -4815
rect 625 -4820 665 -4815
rect 625 -4845 635 -4820
rect 655 -4845 665 -4820
rect 925 -4845 940 -4825
rect 625 -4850 665 -4845
rect 635 -4970 660 -4850
rect 925 -4970 940 -4945
rect 3620 -4950 3635 -4780
rect 3930 -4785 3970 -4780
rect 3930 -4810 3940 -4785
rect 3960 -4810 3970 -4785
rect 4230 -4810 4245 -4790
rect 3930 -4815 3970 -4810
rect 3940 -4935 3965 -4815
rect 4230 -4935 4245 -4910
rect 6925 -4915 6940 -4745
rect 7235 -4750 7275 -4745
rect 7235 -4775 7245 -4750
rect 7265 -4775 7275 -4750
rect 7535 -4775 7550 -4755
rect 7235 -4780 7275 -4775
rect 7245 -4900 7270 -4780
rect 7535 -4900 7550 -4875
rect 10230 -4880 10245 -4710
rect 10540 -4715 10580 -4710
rect 10540 -4740 10550 -4715
rect 10570 -4740 10580 -4715
rect 10840 -4740 10855 -4720
rect 10540 -4745 10580 -4740
rect 10550 -4865 10575 -4745
rect 10840 -4865 10855 -4840
rect 635 -4990 940 -4970
rect 925 -5045 940 -5030
rect 315 -5095 330 -5085
rect 315 -5110 740 -5095
rect 725 -5170 740 -5110
rect 3940 -4955 4245 -4935
rect 4230 -5010 4245 -4995
rect 3620 -5060 3635 -5050
rect 3620 -5075 4045 -5060
rect 925 -5170 940 -5145
rect 4030 -5135 4045 -5075
rect 7245 -4920 7550 -4900
rect 7535 -4975 7550 -4960
rect 6925 -5025 6940 -5015
rect 6925 -5040 7350 -5025
rect 4230 -5135 4245 -5110
rect 7335 -5100 7350 -5040
rect 10550 -4885 10855 -4865
rect 10840 -4940 10855 -4925
rect 10230 -4990 10245 -4980
rect 10230 -5005 10655 -4990
rect 7535 -5100 7550 -5075
rect 10640 -5065 10655 -5005
rect 10840 -5065 10855 -5040
rect 10640 -5080 10855 -5065
rect 7335 -5115 7550 -5100
rect 4030 -5150 4245 -5135
rect 725 -5185 940 -5170
rect 9525 -5510 9540 -5485
rect 6420 -5630 6435 -5605
rect 2975 -5735 2990 -5710
rect 9525 -5980 9540 -5910
rect 9485 -5990 9540 -5980
rect 9485 -6010 9495 -5990
rect 9515 -6010 9540 -5990
rect 9485 -6020 9540 -6010
rect 6420 -6100 6435 -6030
rect 6380 -6110 6435 -6100
rect 9525 -6110 9540 -6020
rect 6380 -6130 6390 -6110
rect 6410 -6130 6435 -6110
rect 2975 -6205 2990 -6135
rect 6380 -6140 6435 -6130
rect 2935 -6215 2990 -6205
rect 2935 -6235 2945 -6215
rect 2965 -6235 2990 -6215
rect 6420 -6230 6435 -6140
rect 2935 -6245 2990 -6235
rect 2975 -6335 2990 -6245
rect 9525 -6335 9540 -6310
rect 6420 -6455 6435 -6430
rect 2975 -6560 2990 -6535
<< polycont >>
rect 130 -2245 160 -2220
rect 1215 -2255 1245 -2230
rect 220 -2405 240 -2380
rect 630 -2410 650 -2390
rect 720 -2490 740 -2470
rect 3435 -2210 3465 -2185
rect 1305 -2415 1325 -2390
rect 1750 -2395 1780 -2370
rect 2215 -2410 2235 -2390
rect 2880 -2365 2910 -2340
rect 2305 -2490 2325 -2470
rect 4520 -2220 4550 -2195
rect 3525 -2370 3545 -2345
rect 3935 -2375 3955 -2355
rect 4025 -2455 4045 -2435
rect 6740 -2175 6770 -2150
rect 4610 -2380 4630 -2355
rect 5055 -2360 5085 -2335
rect 5520 -2375 5540 -2355
rect 6185 -2330 6215 -2305
rect 5610 -2455 5630 -2435
rect 7825 -2185 7855 -2160
rect 6830 -2335 6850 -2310
rect 7240 -2340 7260 -2320
rect 7330 -2420 7350 -2400
rect 10045 -2140 10075 -2115
rect 7915 -2345 7935 -2320
rect 8360 -2325 8390 -2300
rect 8825 -2340 8845 -2320
rect 9490 -2295 9520 -2270
rect 8915 -2420 8935 -2400
rect 11130 -2150 11160 -2125
rect 10135 -2300 10155 -2275
rect 10545 -2305 10565 -2285
rect 10635 -2385 10655 -2365
rect 11220 -2310 11240 -2285
rect 11665 -2290 11695 -2265
rect 12130 -2305 12150 -2285
rect 12795 -2260 12825 -2235
rect 12220 -2385 12240 -2365
rect 315 -3545 345 -3520
rect 685 -3585 705 -3560
rect 3620 -3510 3650 -3485
rect 1840 -4045 1870 -4020
rect 3990 -3550 4010 -3525
rect 6925 -3475 6955 -3450
rect 2210 -4085 2230 -4060
rect 5145 -4010 5175 -3985
rect 7295 -3515 7315 -3490
rect 10230 -3440 10260 -3415
rect 5515 -4050 5535 -4025
rect 2870 -4415 2890 -4395
rect 265 -4805 295 -4780
rect 8450 -3975 8480 -3950
rect 10600 -3480 10620 -3455
rect 8820 -4015 8840 -3990
rect 6200 -4380 6220 -4360
rect 3570 -4770 3600 -4745
rect 11755 -3940 11785 -3915
rect 13785 -3770 13805 -3750
rect 13355 -3810 13375 -3790
rect 12125 -3980 12145 -3955
rect 9515 -4345 9535 -4325
rect 6875 -4735 6905 -4710
rect 10180 -4700 10210 -4675
rect 635 -4845 655 -4820
rect 3940 -4810 3960 -4785
rect 7245 -4775 7265 -4750
rect 10550 -4740 10570 -4715
rect 9495 -6010 9515 -5990
rect 6390 -6130 6410 -6110
rect 2945 -6235 2965 -6215
<< locali >>
rect 12595 -1655 12645 -1640
rect 9290 -1690 9340 -1675
rect 5985 -1725 6035 -1710
rect 2680 -1760 2730 -1745
rect 1550 -1790 1600 -1775
rect 1550 -1815 1565 -1790
rect 1585 -1815 1600 -1790
rect 2680 -1785 2695 -1760
rect 2715 -1785 2730 -1760
rect 2680 -1795 2730 -1785
rect 4855 -1755 4905 -1740
rect 4855 -1780 4870 -1755
rect 4890 -1780 4905 -1755
rect 5985 -1750 6000 -1725
rect 6020 -1750 6035 -1725
rect 5985 -1760 6035 -1750
rect 8160 -1720 8210 -1705
rect 8160 -1745 8175 -1720
rect 8195 -1745 8210 -1720
rect 9290 -1715 9305 -1690
rect 9325 -1715 9340 -1690
rect 9290 -1725 9340 -1715
rect 11465 -1685 11515 -1670
rect 11465 -1710 11480 -1685
rect 11500 -1710 11515 -1685
rect 12595 -1680 12610 -1655
rect 12630 -1680 12645 -1655
rect 12595 -1690 12645 -1680
rect 11465 -1720 11515 -1710
rect 12765 -1725 12950 -1715
rect 12765 -1745 12845 -1725
rect 12865 -1745 12950 -1725
rect 8160 -1755 8210 -1745
rect 9460 -1760 9645 -1750
rect 9460 -1780 9540 -1760
rect 9560 -1780 9645 -1760
rect 4855 -1790 4905 -1780
rect 6155 -1795 6340 -1785
rect 6155 -1815 6235 -1795
rect 6255 -1815 6340 -1795
rect 1550 -1825 1600 -1815
rect 2850 -1830 3035 -1820
rect 2850 -1850 2930 -1830
rect 2950 -1850 3035 -1830
rect -95 -1860 -55 -1850
rect -95 -1885 -85 -1860
rect -65 -1885 -55 -1860
rect -95 -1890 -55 -1885
rect 95 -1860 340 -1850
rect 95 -1885 195 -1860
rect 240 -1885 340 -1860
rect 610 -1865 770 -1855
rect 1720 -1860 1905 -1850
rect 95 -1895 340 -1885
rect 495 -1875 535 -1865
rect 495 -1895 505 -1875
rect 525 -1895 535 -1875
rect 120 -2010 160 -1895
rect 120 -2120 130 -2010
rect 155 -2120 160 -2010
rect 120 -2165 160 -2120
rect 200 -2010 240 -1965
rect 200 -2120 205 -2010
rect 230 -2120 240 -2010
rect 200 -2205 240 -2120
rect 280 -2010 320 -1895
rect 495 -1905 535 -1895
rect 610 -1900 665 -1865
rect 750 -1900 770 -1865
rect 990 -1870 1030 -1860
rect 990 -1895 1000 -1870
rect 1020 -1895 1030 -1870
rect 990 -1900 1030 -1895
rect 1180 -1870 1425 -1860
rect 1180 -1895 1280 -1870
rect 1325 -1895 1425 -1870
rect 280 -2120 285 -2010
rect 310 -2120 320 -2010
rect 280 -2165 320 -2120
rect 610 -1910 770 -1900
rect 1180 -1905 1425 -1895
rect 1720 -1880 1800 -1860
rect 1820 -1880 1905 -1860
rect 2195 -1865 2355 -1855
rect 1720 -1890 1905 -1880
rect 2080 -1875 2120 -1865
rect 610 -1915 655 -1910
rect 610 -2020 650 -1915
rect 80 -2220 170 -2210
rect 80 -2245 130 -2220
rect 160 -2245 170 -2220
rect 80 -2255 170 -2245
rect 200 -2255 320 -2205
rect 280 -2350 320 -2255
rect 610 -2220 615 -2020
rect 645 -2220 650 -2020
rect 610 -2350 650 -2220
rect 770 -2015 810 -1950
rect 770 -2215 775 -2015
rect 805 -2215 810 -2015
rect 1205 -2020 1245 -1905
rect 1205 -2130 1215 -2020
rect 1240 -2130 1245 -2020
rect 1205 -2175 1245 -2130
rect 1285 -2020 1325 -1975
rect 1285 -2130 1290 -2020
rect 1315 -2130 1325 -2020
rect 280 -2360 395 -2350
rect 120 -2380 250 -2370
rect 120 -2405 220 -2380
rect 240 -2405 250 -2380
rect 120 -2415 250 -2405
rect 280 -2380 365 -2360
rect 385 -2380 395 -2360
rect 280 -2390 395 -2380
rect 620 -2390 660 -2385
rect 120 -2505 160 -2465
rect 120 -2615 125 -2505
rect 150 -2615 160 -2505
rect 120 -2685 160 -2615
rect 280 -2500 320 -2390
rect 620 -2410 630 -2390
rect 650 -2410 660 -2390
rect 620 -2415 660 -2410
rect 770 -2445 810 -2215
rect 1285 -2215 1325 -2130
rect 1365 -2020 1405 -1905
rect 1365 -2130 1370 -2020
rect 1395 -2130 1405 -2020
rect 1365 -2175 1405 -2130
rect 1720 -2045 1775 -1890
rect 2080 -1895 2090 -1875
rect 2110 -1895 2120 -1875
rect 2080 -1905 2120 -1895
rect 2195 -1900 2250 -1865
rect 2335 -1900 2355 -1865
rect 2195 -1910 2355 -1900
rect 2850 -1860 3035 -1850
rect 3210 -1825 3250 -1815
rect 3210 -1850 3220 -1825
rect 3240 -1850 3250 -1825
rect 3210 -1855 3250 -1850
rect 3400 -1825 3645 -1815
rect 3400 -1850 3500 -1825
rect 3545 -1850 3645 -1825
rect 3915 -1830 4075 -1820
rect 5025 -1825 5210 -1815
rect 3400 -1860 3645 -1850
rect 3800 -1840 3840 -1830
rect 3800 -1860 3810 -1840
rect 3830 -1860 3840 -1840
rect 2195 -1915 2240 -1910
rect 1720 -2115 1730 -2045
rect 1760 -2115 1775 -2045
rect 1720 -2165 1775 -2115
rect 1835 -2045 1890 -1990
rect 1835 -2115 1850 -2045
rect 1880 -2115 1890 -2045
rect 1205 -2230 1255 -2220
rect 1205 -2255 1215 -2230
rect 1245 -2255 1255 -2230
rect 1205 -2265 1255 -2255
rect 1285 -2265 1405 -2215
rect 1365 -2360 1405 -2265
rect 1365 -2370 1800 -2360
rect 1295 -2390 1335 -2380
rect 1295 -2415 1305 -2390
rect 1325 -2415 1335 -2390
rect 1295 -2425 1335 -2415
rect 1365 -2395 1750 -2370
rect 1780 -2395 1800 -2370
rect 1365 -2400 1800 -2395
rect 1835 -2370 1890 -2115
rect 2195 -2020 2235 -1915
rect 2195 -2220 2200 -2020
rect 2230 -2220 2235 -2020
rect 2195 -2350 2235 -2220
rect 2355 -2015 2395 -1950
rect 2355 -2215 2360 -2015
rect 2390 -2215 2395 -2015
rect 2850 -2015 2905 -1860
rect 2850 -2085 2860 -2015
rect 2890 -2085 2905 -2015
rect 2850 -2135 2905 -2085
rect 2965 -2015 3020 -1960
rect 2965 -2085 2980 -2015
rect 3010 -2085 3020 -2015
rect 1835 -2390 1855 -2370
rect 1875 -2390 1890 -2370
rect 770 -2455 865 -2445
rect 710 -2470 750 -2465
rect 710 -2490 720 -2470
rect 740 -2490 750 -2470
rect 710 -2495 750 -2490
rect 770 -2475 835 -2455
rect 855 -2475 865 -2455
rect 770 -2485 865 -2475
rect 280 -2610 290 -2500
rect 315 -2610 320 -2500
rect 770 -2525 810 -2485
rect 690 -2560 810 -2525
rect 1205 -2515 1245 -2475
rect 280 -2665 320 -2610
rect 610 -2595 650 -2575
rect 610 -2655 615 -2595
rect 640 -2655 650 -2595
rect -55 -2720 160 -2685
rect 610 -2695 650 -2655
rect 690 -2595 730 -2560
rect 690 -2655 700 -2595
rect 725 -2655 730 -2595
rect 690 -2675 730 -2655
rect 770 -2595 810 -2585
rect 770 -2655 775 -2595
rect 800 -2655 810 -2595
rect 770 -2695 810 -2655
rect 1205 -2625 1210 -2515
rect 1235 -2625 1245 -2515
rect 1205 -2695 1245 -2625
rect 1365 -2510 1405 -2400
rect 1365 -2620 1375 -2510
rect 1400 -2620 1405 -2510
rect 1365 -2675 1405 -2620
rect 1725 -2590 1775 -2580
rect 1725 -2660 1735 -2590
rect 1765 -2660 1775 -2590
rect 600 -2700 810 -2695
rect 480 -2710 810 -2700
rect -55 -2730 -15 -2720
rect -55 -2755 -45 -2730
rect -25 -2755 -15 -2730
rect -55 -2760 -15 -2755
rect 120 -2730 320 -2720
rect 120 -2755 185 -2730
rect 235 -2755 320 -2730
rect 480 -2740 490 -2710
rect 535 -2740 680 -2710
rect 480 -2750 680 -2740
rect 740 -2750 810 -2710
rect 600 -2755 810 -2750
rect 1030 -2730 1245 -2695
rect 1725 -2700 1775 -2660
rect 1835 -2590 1890 -2390
rect 2205 -2390 2245 -2385
rect 2205 -2410 2215 -2390
rect 2235 -2410 2245 -2390
rect 2205 -2415 2245 -2410
rect 2355 -2450 2395 -2215
rect 2440 -2340 2930 -2330
rect 2440 -2365 2880 -2340
rect 2910 -2365 2930 -2340
rect 2440 -2370 2930 -2365
rect 2965 -2340 3020 -2085
rect 3425 -1975 3465 -1860
rect 3425 -2085 3435 -1975
rect 3460 -2085 3465 -1975
rect 3425 -2130 3465 -2085
rect 3505 -1975 3545 -1930
rect 3505 -2085 3510 -1975
rect 3535 -2085 3545 -1975
rect 3505 -2170 3545 -2085
rect 3585 -1975 3625 -1860
rect 3800 -1870 3840 -1860
rect 3915 -1865 3970 -1830
rect 4055 -1865 4075 -1830
rect 4295 -1835 4335 -1825
rect 4295 -1860 4305 -1835
rect 4325 -1860 4335 -1835
rect 4295 -1865 4335 -1860
rect 4485 -1835 4730 -1825
rect 4485 -1860 4585 -1835
rect 4630 -1860 4730 -1835
rect 3585 -2085 3590 -1975
rect 3615 -2085 3625 -1975
rect 3585 -2130 3625 -2085
rect 3915 -1875 4075 -1865
rect 4485 -1870 4730 -1860
rect 5025 -1845 5105 -1825
rect 5125 -1845 5210 -1825
rect 5500 -1830 5660 -1820
rect 5025 -1855 5210 -1845
rect 5385 -1840 5425 -1830
rect 3915 -1880 3960 -1875
rect 3915 -1985 3955 -1880
rect 3385 -2185 3475 -2175
rect 3385 -2210 3435 -2185
rect 3465 -2210 3475 -2185
rect 3385 -2220 3475 -2210
rect 3505 -2220 3625 -2170
rect 3585 -2315 3625 -2220
rect 3915 -2185 3920 -1985
rect 3950 -2185 3955 -1985
rect 3915 -2315 3955 -2185
rect 4075 -1980 4115 -1915
rect 4075 -2180 4080 -1980
rect 4110 -2180 4115 -1980
rect 4510 -1985 4550 -1870
rect 4510 -2095 4520 -1985
rect 4545 -2095 4550 -1985
rect 4510 -2140 4550 -2095
rect 4590 -1985 4630 -1940
rect 4590 -2095 4595 -1985
rect 4620 -2095 4630 -1985
rect 3585 -2325 3700 -2315
rect 2965 -2360 2985 -2340
rect 3005 -2360 3020 -2340
rect 2440 -2450 2475 -2370
rect 2295 -2470 2335 -2465
rect 2295 -2490 2305 -2470
rect 2325 -2490 2335 -2470
rect 2295 -2495 2335 -2490
rect 2355 -2485 2475 -2450
rect 2355 -2525 2395 -2485
rect 2275 -2560 2395 -2525
rect 2855 -2560 2905 -2550
rect 1835 -2660 1845 -2590
rect 1875 -2660 1890 -2590
rect 1835 -2670 1890 -2660
rect 2195 -2595 2235 -2575
rect 2195 -2655 2200 -2595
rect 2225 -2655 2235 -2595
rect 2195 -2695 2235 -2655
rect 2275 -2595 2315 -2560
rect 2275 -2655 2285 -2595
rect 2310 -2655 2315 -2595
rect 2275 -2675 2315 -2655
rect 2355 -2595 2395 -2585
rect 2355 -2655 2360 -2595
rect 2385 -2655 2395 -2595
rect 2355 -2695 2395 -2655
rect 2855 -2630 2865 -2560
rect 2895 -2630 2905 -2560
rect 2855 -2670 2905 -2630
rect 2965 -2560 3020 -2360
rect 3425 -2345 3555 -2335
rect 3425 -2370 3525 -2345
rect 3545 -2370 3555 -2345
rect 3425 -2380 3555 -2370
rect 3585 -2345 3670 -2325
rect 3690 -2345 3700 -2325
rect 3585 -2355 3700 -2345
rect 3925 -2355 3965 -2350
rect 2965 -2630 2975 -2560
rect 3005 -2630 3020 -2560
rect 2965 -2640 3020 -2630
rect 3425 -2470 3465 -2430
rect 3425 -2580 3430 -2470
rect 3455 -2580 3465 -2470
rect 3425 -2650 3465 -2580
rect 3585 -2465 3625 -2355
rect 3925 -2375 3935 -2355
rect 3955 -2375 3965 -2355
rect 3925 -2380 3965 -2375
rect 4075 -2410 4115 -2180
rect 4590 -2180 4630 -2095
rect 4670 -1985 4710 -1870
rect 4670 -2095 4675 -1985
rect 4700 -2095 4710 -1985
rect 4670 -2140 4710 -2095
rect 5025 -2010 5080 -1855
rect 5385 -1860 5395 -1840
rect 5415 -1860 5425 -1840
rect 5385 -1870 5425 -1860
rect 5500 -1865 5555 -1830
rect 5640 -1865 5660 -1830
rect 5500 -1875 5660 -1865
rect 6155 -1825 6340 -1815
rect 6515 -1790 6555 -1780
rect 6515 -1815 6525 -1790
rect 6545 -1815 6555 -1790
rect 6515 -1820 6555 -1815
rect 6705 -1790 6950 -1780
rect 6705 -1815 6805 -1790
rect 6850 -1815 6950 -1790
rect 7220 -1795 7380 -1785
rect 8330 -1790 8515 -1780
rect 6705 -1825 6950 -1815
rect 7105 -1805 7145 -1795
rect 7105 -1825 7115 -1805
rect 7135 -1825 7145 -1805
rect 5500 -1880 5545 -1875
rect 5025 -2080 5035 -2010
rect 5065 -2080 5080 -2010
rect 5025 -2130 5080 -2080
rect 5140 -2010 5195 -1955
rect 5140 -2080 5155 -2010
rect 5185 -2080 5195 -2010
rect 4445 -2195 4560 -2185
rect 4445 -2220 4520 -2195
rect 4550 -2220 4560 -2195
rect 4445 -2230 4560 -2220
rect 4590 -2230 4710 -2180
rect 4670 -2325 4710 -2230
rect 4670 -2335 5105 -2325
rect 4600 -2355 4640 -2345
rect 4600 -2380 4610 -2355
rect 4630 -2380 4640 -2355
rect 4600 -2390 4640 -2380
rect 4670 -2360 5055 -2335
rect 5085 -2360 5105 -2335
rect 4670 -2365 5105 -2360
rect 5140 -2335 5195 -2080
rect 5500 -1985 5540 -1880
rect 5500 -2185 5505 -1985
rect 5535 -2185 5540 -1985
rect 5500 -2315 5540 -2185
rect 5660 -1980 5700 -1915
rect 5660 -2180 5665 -1980
rect 5695 -2180 5700 -1980
rect 6155 -1980 6210 -1825
rect 6155 -2050 6165 -1980
rect 6195 -2050 6210 -1980
rect 6155 -2100 6210 -2050
rect 6270 -1980 6325 -1925
rect 6270 -2050 6285 -1980
rect 6315 -2050 6325 -1980
rect 5140 -2355 5160 -2335
rect 5180 -2355 5195 -2335
rect 4075 -2420 4170 -2410
rect 4015 -2435 4055 -2430
rect 4015 -2455 4025 -2435
rect 4045 -2455 4055 -2435
rect 4015 -2460 4055 -2455
rect 4075 -2440 4140 -2420
rect 4160 -2440 4170 -2420
rect 4075 -2450 4170 -2440
rect 3585 -2575 3595 -2465
rect 3620 -2575 3625 -2465
rect 4075 -2490 4115 -2450
rect 3995 -2525 4115 -2490
rect 4510 -2480 4550 -2440
rect 3585 -2630 3625 -2575
rect 3915 -2560 3955 -2540
rect 3915 -2620 3920 -2560
rect 3945 -2620 3955 -2560
rect 2185 -2700 2395 -2695
rect 1570 -2715 1775 -2700
rect 2065 -2710 2395 -2700
rect 1570 -2725 1905 -2715
rect 1030 -2740 1070 -2730
rect 120 -2765 320 -2755
rect 1030 -2765 1040 -2740
rect 1060 -2765 1070 -2740
rect 1030 -2770 1070 -2765
rect 1205 -2740 1405 -2730
rect 1205 -2765 1270 -2740
rect 1320 -2765 1405 -2740
rect 1205 -2775 1405 -2765
rect 1570 -2735 1795 -2725
rect 1570 -2740 1610 -2735
rect 1570 -2765 1580 -2740
rect 1600 -2765 1610 -2740
rect 1725 -2745 1795 -2735
rect 1820 -2745 1905 -2725
rect 1725 -2750 1905 -2745
rect 2065 -2740 2075 -2710
rect 2120 -2740 2265 -2710
rect 2065 -2750 2265 -2740
rect 2325 -2750 2395 -2710
rect 2700 -2685 2905 -2670
rect 3250 -2685 3465 -2650
rect 3915 -2660 3955 -2620
rect 3995 -2560 4035 -2525
rect 3995 -2620 4005 -2560
rect 4030 -2620 4035 -2560
rect 3995 -2640 4035 -2620
rect 4075 -2560 4115 -2550
rect 4075 -2620 4080 -2560
rect 4105 -2620 4115 -2560
rect 4075 -2660 4115 -2620
rect 4510 -2590 4515 -2480
rect 4540 -2590 4550 -2480
rect 4510 -2660 4550 -2590
rect 4670 -2475 4710 -2365
rect 4670 -2585 4680 -2475
rect 4705 -2585 4710 -2475
rect 4670 -2640 4710 -2585
rect 5030 -2555 5080 -2545
rect 5030 -2625 5040 -2555
rect 5070 -2625 5080 -2555
rect 3905 -2665 4115 -2660
rect 3785 -2675 4115 -2665
rect 2700 -2695 3035 -2685
rect 2700 -2705 2925 -2695
rect 2700 -2710 2740 -2705
rect 2700 -2735 2710 -2710
rect 2730 -2735 2740 -2710
rect 2855 -2715 2925 -2705
rect 2950 -2715 3035 -2695
rect 2855 -2720 3035 -2715
rect 3250 -2695 3290 -2685
rect 3250 -2720 3260 -2695
rect 3280 -2720 3290 -2695
rect 3250 -2725 3290 -2720
rect 3425 -2695 3625 -2685
rect 3425 -2720 3490 -2695
rect 3540 -2720 3625 -2695
rect 3785 -2705 3795 -2675
rect 3840 -2705 3985 -2675
rect 3785 -2715 3985 -2705
rect 4045 -2715 4115 -2675
rect 3905 -2720 4115 -2715
rect 4335 -2695 4550 -2660
rect 5030 -2665 5080 -2625
rect 5140 -2555 5195 -2355
rect 5510 -2355 5550 -2350
rect 5510 -2375 5520 -2355
rect 5540 -2375 5550 -2355
rect 5510 -2380 5550 -2375
rect 5660 -2415 5700 -2180
rect 5745 -2305 6235 -2295
rect 5745 -2330 6185 -2305
rect 6215 -2330 6235 -2305
rect 5745 -2335 6235 -2330
rect 6270 -2305 6325 -2050
rect 6730 -1940 6770 -1825
rect 6730 -2050 6740 -1940
rect 6765 -2050 6770 -1940
rect 6730 -2095 6770 -2050
rect 6810 -1940 6850 -1895
rect 6810 -2050 6815 -1940
rect 6840 -2050 6850 -1940
rect 6810 -2135 6850 -2050
rect 6890 -1940 6930 -1825
rect 7105 -1835 7145 -1825
rect 7220 -1830 7275 -1795
rect 7360 -1830 7380 -1795
rect 7600 -1800 7640 -1790
rect 7600 -1825 7610 -1800
rect 7630 -1825 7640 -1800
rect 7600 -1830 7640 -1825
rect 7790 -1800 8035 -1790
rect 7790 -1825 7890 -1800
rect 7935 -1825 8035 -1800
rect 6890 -2050 6895 -1940
rect 6920 -2050 6930 -1940
rect 6890 -2095 6930 -2050
rect 7220 -1840 7380 -1830
rect 7790 -1835 8035 -1825
rect 8330 -1810 8410 -1790
rect 8430 -1810 8515 -1790
rect 8805 -1795 8965 -1785
rect 8330 -1820 8515 -1810
rect 8690 -1805 8730 -1795
rect 7220 -1845 7265 -1840
rect 7220 -1950 7260 -1845
rect 6690 -2150 6780 -2140
rect 6690 -2175 6740 -2150
rect 6770 -2175 6780 -2150
rect 6690 -2185 6780 -2175
rect 6810 -2185 6930 -2135
rect 6890 -2280 6930 -2185
rect 7220 -2150 7225 -1950
rect 7255 -2150 7260 -1950
rect 7220 -2280 7260 -2150
rect 7380 -1945 7420 -1880
rect 7380 -2145 7385 -1945
rect 7415 -2145 7420 -1945
rect 7815 -1950 7855 -1835
rect 7815 -2060 7825 -1950
rect 7850 -2060 7855 -1950
rect 7815 -2105 7855 -2060
rect 7895 -1950 7935 -1905
rect 7895 -2060 7900 -1950
rect 7925 -2060 7935 -1950
rect 6890 -2290 7005 -2280
rect 6270 -2325 6290 -2305
rect 6310 -2325 6325 -2305
rect 5745 -2415 5780 -2335
rect 5600 -2435 5640 -2430
rect 5600 -2455 5610 -2435
rect 5630 -2455 5640 -2435
rect 5600 -2460 5640 -2455
rect 5660 -2450 5780 -2415
rect 5660 -2490 5700 -2450
rect 5580 -2525 5700 -2490
rect 6160 -2525 6210 -2515
rect 5140 -2625 5150 -2555
rect 5180 -2625 5195 -2555
rect 5140 -2635 5195 -2625
rect 5500 -2560 5540 -2540
rect 5500 -2620 5505 -2560
rect 5530 -2620 5540 -2560
rect 5500 -2660 5540 -2620
rect 5580 -2560 5620 -2525
rect 5580 -2620 5590 -2560
rect 5615 -2620 5620 -2560
rect 5580 -2640 5620 -2620
rect 5660 -2560 5700 -2550
rect 5660 -2620 5665 -2560
rect 5690 -2620 5700 -2560
rect 5660 -2660 5700 -2620
rect 6160 -2595 6170 -2525
rect 6200 -2595 6210 -2525
rect 6160 -2635 6210 -2595
rect 6270 -2525 6325 -2325
rect 6730 -2310 6860 -2300
rect 6730 -2335 6830 -2310
rect 6850 -2335 6860 -2310
rect 6730 -2345 6860 -2335
rect 6890 -2310 6975 -2290
rect 6995 -2310 7005 -2290
rect 6890 -2320 7005 -2310
rect 7230 -2320 7270 -2315
rect 6270 -2595 6280 -2525
rect 6310 -2595 6325 -2525
rect 6270 -2605 6325 -2595
rect 6730 -2435 6770 -2395
rect 6730 -2545 6735 -2435
rect 6760 -2545 6770 -2435
rect 6730 -2615 6770 -2545
rect 6890 -2430 6930 -2320
rect 7230 -2340 7240 -2320
rect 7260 -2340 7270 -2320
rect 7230 -2345 7270 -2340
rect 7380 -2375 7420 -2145
rect 7895 -2145 7935 -2060
rect 7975 -1950 8015 -1835
rect 7975 -2060 7980 -1950
rect 8005 -2060 8015 -1950
rect 7975 -2105 8015 -2060
rect 8330 -1975 8385 -1820
rect 8690 -1825 8700 -1805
rect 8720 -1825 8730 -1805
rect 8690 -1835 8730 -1825
rect 8805 -1830 8860 -1795
rect 8945 -1830 8965 -1795
rect 8805 -1840 8965 -1830
rect 9460 -1790 9645 -1780
rect 9820 -1755 9860 -1745
rect 9820 -1780 9830 -1755
rect 9850 -1780 9860 -1755
rect 9820 -1785 9860 -1780
rect 10010 -1755 10255 -1745
rect 10010 -1780 10110 -1755
rect 10155 -1780 10255 -1755
rect 10525 -1760 10685 -1750
rect 11635 -1755 11820 -1745
rect 10010 -1790 10255 -1780
rect 10410 -1770 10450 -1760
rect 10410 -1790 10420 -1770
rect 10440 -1790 10450 -1770
rect 8805 -1845 8850 -1840
rect 8330 -2045 8340 -1975
rect 8370 -2045 8385 -1975
rect 8330 -2095 8385 -2045
rect 8445 -1975 8500 -1920
rect 8445 -2045 8460 -1975
rect 8490 -2045 8500 -1975
rect 7750 -2160 7865 -2150
rect 7750 -2185 7825 -2160
rect 7855 -2185 7865 -2160
rect 7750 -2195 7865 -2185
rect 7895 -2195 8015 -2145
rect 7975 -2290 8015 -2195
rect 7975 -2300 8410 -2290
rect 7905 -2320 7945 -2310
rect 7905 -2345 7915 -2320
rect 7935 -2345 7945 -2320
rect 7905 -2355 7945 -2345
rect 7975 -2325 8360 -2300
rect 8390 -2325 8410 -2300
rect 7975 -2330 8410 -2325
rect 8445 -2300 8500 -2045
rect 8805 -1950 8845 -1845
rect 8805 -2150 8810 -1950
rect 8840 -2150 8845 -1950
rect 8805 -2280 8845 -2150
rect 8965 -1945 9005 -1880
rect 8965 -2145 8970 -1945
rect 9000 -2145 9005 -1945
rect 9460 -1945 9515 -1790
rect 9460 -2015 9470 -1945
rect 9500 -2015 9515 -1945
rect 9460 -2065 9515 -2015
rect 9575 -1945 9630 -1890
rect 9575 -2015 9590 -1945
rect 9620 -2015 9630 -1945
rect 8445 -2320 8465 -2300
rect 8485 -2320 8500 -2300
rect 7380 -2385 7475 -2375
rect 7320 -2400 7360 -2395
rect 7320 -2420 7330 -2400
rect 7350 -2420 7360 -2400
rect 7320 -2425 7360 -2420
rect 7380 -2405 7445 -2385
rect 7465 -2405 7475 -2385
rect 7380 -2415 7475 -2405
rect 6890 -2540 6900 -2430
rect 6925 -2540 6930 -2430
rect 7380 -2455 7420 -2415
rect 7300 -2490 7420 -2455
rect 7815 -2445 7855 -2405
rect 6890 -2595 6930 -2540
rect 7220 -2525 7260 -2505
rect 7220 -2585 7225 -2525
rect 7250 -2585 7260 -2525
rect 5490 -2665 5700 -2660
rect 4875 -2680 5080 -2665
rect 5370 -2675 5700 -2665
rect 4875 -2690 5210 -2680
rect 4335 -2705 4375 -2695
rect 3425 -2730 3625 -2720
rect 4335 -2730 4345 -2705
rect 4365 -2730 4375 -2705
rect 4335 -2735 4375 -2730
rect 4510 -2705 4710 -2695
rect 4510 -2730 4575 -2705
rect 4625 -2730 4710 -2705
rect 2700 -2740 2740 -2735
rect 4510 -2740 4710 -2730
rect 4875 -2700 5100 -2690
rect 4875 -2705 4915 -2700
rect 4875 -2730 4885 -2705
rect 4905 -2730 4915 -2705
rect 5030 -2710 5100 -2700
rect 5125 -2710 5210 -2690
rect 5030 -2715 5210 -2710
rect 5370 -2705 5380 -2675
rect 5425 -2705 5570 -2675
rect 5370 -2715 5570 -2705
rect 5630 -2715 5700 -2675
rect 6005 -2650 6210 -2635
rect 6555 -2650 6770 -2615
rect 7220 -2625 7260 -2585
rect 7300 -2525 7340 -2490
rect 7300 -2585 7310 -2525
rect 7335 -2585 7340 -2525
rect 7300 -2605 7340 -2585
rect 7380 -2525 7420 -2515
rect 7380 -2585 7385 -2525
rect 7410 -2585 7420 -2525
rect 7380 -2625 7420 -2585
rect 7815 -2555 7820 -2445
rect 7845 -2555 7855 -2445
rect 7815 -2625 7855 -2555
rect 7975 -2440 8015 -2330
rect 7975 -2550 7985 -2440
rect 8010 -2550 8015 -2440
rect 7975 -2605 8015 -2550
rect 8335 -2520 8385 -2510
rect 8335 -2590 8345 -2520
rect 8375 -2590 8385 -2520
rect 7210 -2630 7420 -2625
rect 7090 -2640 7420 -2630
rect 6005 -2660 6340 -2650
rect 6005 -2670 6230 -2660
rect 6005 -2675 6045 -2670
rect 6005 -2700 6015 -2675
rect 6035 -2700 6045 -2675
rect 6160 -2680 6230 -2670
rect 6255 -2680 6340 -2660
rect 6160 -2685 6340 -2680
rect 6555 -2660 6595 -2650
rect 6555 -2685 6565 -2660
rect 6585 -2685 6595 -2660
rect 6555 -2690 6595 -2685
rect 6730 -2660 6930 -2650
rect 6730 -2685 6795 -2660
rect 6845 -2685 6930 -2660
rect 7090 -2670 7100 -2640
rect 7145 -2670 7290 -2640
rect 7090 -2680 7290 -2670
rect 7350 -2680 7420 -2640
rect 7210 -2685 7420 -2680
rect 7640 -2660 7855 -2625
rect 8335 -2630 8385 -2590
rect 8445 -2520 8500 -2320
rect 8815 -2320 8855 -2315
rect 8815 -2340 8825 -2320
rect 8845 -2340 8855 -2320
rect 8815 -2345 8855 -2340
rect 8965 -2380 9005 -2145
rect 9050 -2270 9540 -2260
rect 9050 -2295 9490 -2270
rect 9520 -2295 9540 -2270
rect 9050 -2300 9540 -2295
rect 9575 -2270 9630 -2015
rect 10035 -1905 10075 -1790
rect 10035 -2015 10045 -1905
rect 10070 -2015 10075 -1905
rect 10035 -2060 10075 -2015
rect 10115 -1905 10155 -1860
rect 10115 -2015 10120 -1905
rect 10145 -2015 10155 -1905
rect 10115 -2100 10155 -2015
rect 10195 -1905 10235 -1790
rect 10410 -1800 10450 -1790
rect 10525 -1795 10580 -1760
rect 10665 -1795 10685 -1760
rect 10905 -1765 10945 -1755
rect 10905 -1790 10915 -1765
rect 10935 -1790 10945 -1765
rect 10905 -1795 10945 -1790
rect 11095 -1765 11340 -1755
rect 11095 -1790 11195 -1765
rect 11240 -1790 11340 -1765
rect 10195 -2015 10200 -1905
rect 10225 -2015 10235 -1905
rect 10195 -2060 10235 -2015
rect 10525 -1805 10685 -1795
rect 11095 -1800 11340 -1790
rect 11635 -1775 11715 -1755
rect 11735 -1775 11820 -1755
rect 12110 -1760 12270 -1750
rect 11635 -1785 11820 -1775
rect 11995 -1770 12035 -1760
rect 10525 -1810 10570 -1805
rect 10525 -1915 10565 -1810
rect 9995 -2115 10085 -2105
rect 9995 -2140 10045 -2115
rect 10075 -2140 10085 -2115
rect 9995 -2150 10085 -2140
rect 10115 -2150 10235 -2100
rect 10195 -2245 10235 -2150
rect 10525 -2115 10530 -1915
rect 10560 -2115 10565 -1915
rect 10525 -2245 10565 -2115
rect 10685 -1910 10725 -1845
rect 10685 -2110 10690 -1910
rect 10720 -2110 10725 -1910
rect 11120 -1915 11160 -1800
rect 11120 -2025 11130 -1915
rect 11155 -2025 11160 -1915
rect 11120 -2070 11160 -2025
rect 11200 -1915 11240 -1870
rect 11200 -2025 11205 -1915
rect 11230 -2025 11240 -1915
rect 10195 -2255 10310 -2245
rect 9575 -2290 9595 -2270
rect 9615 -2290 9630 -2270
rect 9050 -2380 9085 -2300
rect 8905 -2400 8945 -2395
rect 8905 -2420 8915 -2400
rect 8935 -2420 8945 -2400
rect 8905 -2425 8945 -2420
rect 8965 -2415 9085 -2380
rect 8965 -2455 9005 -2415
rect 8885 -2490 9005 -2455
rect 9465 -2490 9515 -2480
rect 8445 -2590 8455 -2520
rect 8485 -2590 8500 -2520
rect 8445 -2600 8500 -2590
rect 8805 -2525 8845 -2505
rect 8805 -2585 8810 -2525
rect 8835 -2585 8845 -2525
rect 8805 -2625 8845 -2585
rect 8885 -2525 8925 -2490
rect 8885 -2585 8895 -2525
rect 8920 -2585 8925 -2525
rect 8885 -2605 8925 -2585
rect 8965 -2525 9005 -2515
rect 8965 -2585 8970 -2525
rect 8995 -2585 9005 -2525
rect 8965 -2625 9005 -2585
rect 9465 -2560 9475 -2490
rect 9505 -2560 9515 -2490
rect 9465 -2600 9515 -2560
rect 9575 -2490 9630 -2290
rect 10035 -2275 10165 -2265
rect 10035 -2300 10135 -2275
rect 10155 -2300 10165 -2275
rect 10035 -2310 10165 -2300
rect 10195 -2275 10280 -2255
rect 10300 -2275 10310 -2255
rect 10195 -2285 10310 -2275
rect 10535 -2285 10575 -2280
rect 9575 -2560 9585 -2490
rect 9615 -2560 9630 -2490
rect 9575 -2570 9630 -2560
rect 10035 -2400 10075 -2360
rect 10035 -2510 10040 -2400
rect 10065 -2510 10075 -2400
rect 10035 -2580 10075 -2510
rect 10195 -2395 10235 -2285
rect 10535 -2305 10545 -2285
rect 10565 -2305 10575 -2285
rect 10535 -2310 10575 -2305
rect 10685 -2340 10725 -2110
rect 11200 -2110 11240 -2025
rect 11280 -1915 11320 -1800
rect 11280 -2025 11285 -1915
rect 11310 -2025 11320 -1915
rect 11280 -2070 11320 -2025
rect 11635 -1940 11690 -1785
rect 11995 -1790 12005 -1770
rect 12025 -1790 12035 -1770
rect 11995 -1800 12035 -1790
rect 12110 -1795 12165 -1760
rect 12250 -1795 12270 -1760
rect 12110 -1805 12270 -1795
rect 12765 -1755 12950 -1745
rect 12110 -1810 12155 -1805
rect 11635 -2010 11645 -1940
rect 11675 -2010 11690 -1940
rect 11635 -2060 11690 -2010
rect 11750 -1940 11805 -1885
rect 11750 -2010 11765 -1940
rect 11795 -2010 11805 -1940
rect 11055 -2125 11170 -2115
rect 11055 -2150 11130 -2125
rect 11160 -2150 11170 -2125
rect 11055 -2160 11170 -2150
rect 11200 -2160 11320 -2110
rect 11280 -2255 11320 -2160
rect 11280 -2265 11715 -2255
rect 11210 -2285 11250 -2275
rect 11210 -2310 11220 -2285
rect 11240 -2310 11250 -2285
rect 11210 -2320 11250 -2310
rect 11280 -2290 11665 -2265
rect 11695 -2290 11715 -2265
rect 11280 -2295 11715 -2290
rect 11750 -2265 11805 -2010
rect 12110 -1915 12150 -1810
rect 12110 -2115 12115 -1915
rect 12145 -2115 12150 -1915
rect 12110 -2245 12150 -2115
rect 12270 -1910 12310 -1845
rect 12270 -2110 12275 -1910
rect 12305 -2110 12310 -1910
rect 12765 -1910 12820 -1755
rect 12765 -1980 12775 -1910
rect 12805 -1980 12820 -1910
rect 12765 -2030 12820 -1980
rect 12880 -1910 12935 -1855
rect 12880 -1980 12895 -1910
rect 12925 -1980 12935 -1910
rect 11750 -2285 11770 -2265
rect 11790 -2285 11805 -2265
rect 10685 -2350 10780 -2340
rect 10625 -2365 10665 -2360
rect 10625 -2385 10635 -2365
rect 10655 -2385 10665 -2365
rect 10625 -2390 10665 -2385
rect 10685 -2370 10750 -2350
rect 10770 -2370 10780 -2350
rect 10685 -2380 10780 -2370
rect 10195 -2505 10205 -2395
rect 10230 -2505 10235 -2395
rect 10685 -2420 10725 -2380
rect 10605 -2455 10725 -2420
rect 11120 -2410 11160 -2370
rect 10195 -2560 10235 -2505
rect 10525 -2490 10565 -2470
rect 10525 -2550 10530 -2490
rect 10555 -2550 10565 -2490
rect 8795 -2630 9005 -2625
rect 8180 -2645 8385 -2630
rect 8675 -2640 9005 -2630
rect 8180 -2655 8515 -2645
rect 7640 -2670 7680 -2660
rect 6730 -2695 6930 -2685
rect 7640 -2695 7650 -2670
rect 7670 -2695 7680 -2670
rect 7640 -2700 7680 -2695
rect 7815 -2670 8015 -2660
rect 7815 -2695 7880 -2670
rect 7930 -2695 8015 -2670
rect 6005 -2705 6045 -2700
rect 7815 -2705 8015 -2695
rect 8180 -2665 8405 -2655
rect 8180 -2670 8220 -2665
rect 8180 -2695 8190 -2670
rect 8210 -2695 8220 -2670
rect 8335 -2675 8405 -2665
rect 8430 -2675 8515 -2655
rect 8335 -2680 8515 -2675
rect 8675 -2670 8685 -2640
rect 8730 -2670 8875 -2640
rect 8675 -2680 8875 -2670
rect 8935 -2680 9005 -2640
rect 9310 -2615 9515 -2600
rect 9860 -2615 10075 -2580
rect 10525 -2590 10565 -2550
rect 10605 -2490 10645 -2455
rect 10605 -2550 10615 -2490
rect 10640 -2550 10645 -2490
rect 10605 -2570 10645 -2550
rect 10685 -2490 10725 -2480
rect 10685 -2550 10690 -2490
rect 10715 -2550 10725 -2490
rect 10685 -2590 10725 -2550
rect 11120 -2520 11125 -2410
rect 11150 -2520 11160 -2410
rect 11120 -2590 11160 -2520
rect 11280 -2405 11320 -2295
rect 11280 -2515 11290 -2405
rect 11315 -2515 11320 -2405
rect 11280 -2570 11320 -2515
rect 11640 -2485 11690 -2475
rect 11640 -2555 11650 -2485
rect 11680 -2555 11690 -2485
rect 10515 -2595 10725 -2590
rect 10395 -2605 10725 -2595
rect 9310 -2625 9645 -2615
rect 9310 -2635 9535 -2625
rect 9310 -2640 9350 -2635
rect 9310 -2665 9320 -2640
rect 9340 -2665 9350 -2640
rect 9465 -2645 9535 -2635
rect 9560 -2645 9645 -2625
rect 9465 -2650 9645 -2645
rect 9860 -2625 9900 -2615
rect 9860 -2650 9870 -2625
rect 9890 -2650 9900 -2625
rect 9860 -2655 9900 -2650
rect 10035 -2625 10235 -2615
rect 10035 -2650 10100 -2625
rect 10150 -2650 10235 -2625
rect 10395 -2635 10405 -2605
rect 10450 -2635 10595 -2605
rect 10395 -2645 10595 -2635
rect 10655 -2645 10725 -2605
rect 10515 -2650 10725 -2645
rect 10945 -2625 11160 -2590
rect 11640 -2595 11690 -2555
rect 11750 -2485 11805 -2285
rect 12120 -2285 12160 -2280
rect 12120 -2305 12130 -2285
rect 12150 -2305 12160 -2285
rect 12120 -2310 12160 -2305
rect 12270 -2345 12310 -2110
rect 12355 -2235 12845 -2225
rect 12355 -2260 12795 -2235
rect 12825 -2260 12845 -2235
rect 12355 -2265 12845 -2260
rect 12880 -2235 12935 -1980
rect 12880 -2255 12900 -2235
rect 12920 -2255 12935 -2235
rect 12355 -2345 12390 -2265
rect 12210 -2365 12250 -2360
rect 12210 -2385 12220 -2365
rect 12240 -2385 12250 -2365
rect 12210 -2390 12250 -2385
rect 12270 -2380 12390 -2345
rect 12270 -2420 12310 -2380
rect 12190 -2455 12310 -2420
rect 12770 -2455 12820 -2445
rect 11750 -2555 11760 -2485
rect 11790 -2555 11805 -2485
rect 11750 -2565 11805 -2555
rect 12110 -2490 12150 -2470
rect 12110 -2550 12115 -2490
rect 12140 -2550 12150 -2490
rect 12110 -2590 12150 -2550
rect 12190 -2490 12230 -2455
rect 12190 -2550 12200 -2490
rect 12225 -2550 12230 -2490
rect 12190 -2570 12230 -2550
rect 12270 -2490 12310 -2480
rect 12270 -2550 12275 -2490
rect 12300 -2550 12310 -2490
rect 12270 -2590 12310 -2550
rect 12770 -2525 12780 -2455
rect 12810 -2525 12820 -2455
rect 12770 -2565 12820 -2525
rect 12880 -2455 12935 -2255
rect 12880 -2525 12890 -2455
rect 12920 -2525 12935 -2455
rect 12880 -2535 12935 -2525
rect 12100 -2595 12310 -2590
rect 11485 -2610 11690 -2595
rect 11980 -2605 12310 -2595
rect 11485 -2620 11820 -2610
rect 10945 -2635 10985 -2625
rect 10035 -2660 10235 -2650
rect 10945 -2660 10955 -2635
rect 10975 -2660 10985 -2635
rect 10945 -2665 10985 -2660
rect 11120 -2635 11320 -2625
rect 11120 -2660 11185 -2635
rect 11235 -2660 11320 -2635
rect 9310 -2670 9350 -2665
rect 11120 -2670 11320 -2660
rect 11485 -2630 11710 -2620
rect 11485 -2635 11525 -2630
rect 11485 -2660 11495 -2635
rect 11515 -2660 11525 -2635
rect 11640 -2640 11710 -2630
rect 11735 -2640 11820 -2620
rect 11640 -2645 11820 -2640
rect 11980 -2635 11990 -2605
rect 12035 -2635 12180 -2605
rect 11980 -2645 12180 -2635
rect 12240 -2645 12310 -2605
rect 12615 -2580 12820 -2565
rect 12615 -2590 12950 -2580
rect 12615 -2600 12840 -2590
rect 12615 -2605 12655 -2600
rect 12615 -2630 12625 -2605
rect 12645 -2630 12655 -2605
rect 12770 -2610 12840 -2600
rect 12865 -2610 12950 -2590
rect 12770 -2615 12950 -2610
rect 12615 -2635 12655 -2630
rect 12100 -2650 12310 -2645
rect 11485 -2665 11525 -2660
rect 8795 -2685 9005 -2680
rect 8180 -2700 8220 -2695
rect 5490 -2720 5700 -2715
rect 4875 -2735 4915 -2730
rect 2185 -2755 2395 -2750
rect 1570 -2770 1610 -2765
rect 10848 -2810 10898 -2795
rect 7543 -2845 7593 -2830
rect 4238 -2880 4288 -2865
rect 933 -2915 983 -2900
rect 115 -2940 165 -2925
rect 115 -2965 130 -2940
rect 150 -2965 165 -2940
rect 933 -2940 948 -2915
rect 968 -2940 983 -2915
rect 3420 -2905 3470 -2890
rect 3420 -2930 3435 -2905
rect 3455 -2930 3470 -2905
rect 4238 -2905 4253 -2880
rect 4273 -2905 4288 -2880
rect 6725 -2870 6775 -2855
rect 6725 -2895 6740 -2870
rect 6760 -2895 6775 -2870
rect 7543 -2870 7558 -2845
rect 7578 -2870 7593 -2845
rect 10030 -2835 10080 -2820
rect 10030 -2860 10045 -2835
rect 10065 -2860 10080 -2835
rect 10848 -2835 10863 -2810
rect 10883 -2835 10898 -2810
rect 10848 -2845 10898 -2835
rect 10030 -2870 10080 -2860
rect 7543 -2880 7593 -2870
rect 10850 -2895 10890 -2885
rect 6725 -2905 6775 -2895
rect 10200 -2905 10385 -2895
rect 4238 -2915 4288 -2905
rect 7545 -2930 7585 -2920
rect 3420 -2940 3470 -2930
rect 6895 -2940 7080 -2930
rect 933 -2950 983 -2940
rect 4240 -2965 4280 -2955
rect 115 -2975 165 -2965
rect 3590 -2975 3775 -2965
rect 935 -3000 975 -2990
rect 285 -3010 470 -3000
rect 285 -3030 365 -3010
rect 385 -3030 470 -3010
rect 285 -3040 470 -3030
rect 285 -3195 340 -3040
rect 935 -3080 945 -3000
rect 965 -3080 975 -3000
rect 935 -3130 975 -3080
rect 285 -3265 295 -3195
rect 325 -3265 340 -3195
rect 285 -3315 340 -3265
rect 400 -3195 455 -3140
rect 400 -3265 415 -3195
rect 445 -3265 455 -3195
rect 130 -3520 365 -3510
rect 130 -3545 315 -3520
rect 345 -3545 365 -3520
rect 130 -3550 365 -3545
rect 400 -3565 455 -3265
rect 935 -3150 945 -3130
rect 965 -3150 975 -3130
rect 935 -3200 975 -3150
rect 935 -3280 945 -3200
rect 965 -3280 975 -3200
rect 935 -3290 975 -3280
rect 1000 -3000 1035 -2990
rect 1000 -3080 1005 -3000
rect 1025 -3080 1035 -3000
rect 1000 -3200 1035 -3080
rect 1000 -3280 1010 -3200
rect 1030 -3280 1035 -3200
rect 3590 -2995 3670 -2975
rect 3690 -2995 3775 -2975
rect 3590 -3005 3775 -2995
rect 3590 -3160 3645 -3005
rect 4240 -3045 4250 -2965
rect 4270 -3045 4280 -2965
rect 4240 -3095 4280 -3045
rect 3590 -3230 3600 -3160
rect 3630 -3230 3645 -3160
rect 3590 -3280 3645 -3230
rect 3705 -3160 3760 -3105
rect 3705 -3230 3720 -3160
rect 3750 -3230 3760 -3160
rect 1000 -3375 1035 -3280
rect 1450 -3375 2375 -3350
rect 1000 -3380 2375 -3375
rect 1000 -3415 1470 -3380
rect 928 -3510 978 -3495
rect 928 -3535 943 -3510
rect 963 -3535 978 -3510
rect 928 -3545 978 -3535
rect 675 -3560 715 -3555
rect 675 -3565 685 -3560
rect 400 -3585 685 -3565
rect 705 -3585 715 -3560
rect 1000 -3585 1035 -3415
rect 1640 -3440 1690 -3425
rect 1640 -3465 1655 -3440
rect 1675 -3465 1690 -3440
rect 1640 -3475 1690 -3465
rect 290 -3740 340 -3730
rect 290 -3810 300 -3740
rect 330 -3810 340 -3740
rect 290 -3850 340 -3810
rect 400 -3740 455 -3585
rect 675 -3590 715 -3585
rect 400 -3810 410 -3740
rect 440 -3810 455 -3740
rect 400 -3820 455 -3810
rect 930 -3595 970 -3585
rect 930 -3675 940 -3595
rect 960 -3675 970 -3595
rect 930 -3745 970 -3675
rect 930 -3765 940 -3745
rect 960 -3765 970 -3745
rect 930 -3795 970 -3765
rect 135 -3865 340 -3850
rect 135 -3875 470 -3865
rect 135 -3885 360 -3875
rect 135 -3890 175 -3885
rect 135 -3915 145 -3890
rect 165 -3915 175 -3890
rect 290 -3895 360 -3885
rect 385 -3895 470 -3875
rect 930 -3875 940 -3795
rect 960 -3875 970 -3795
rect 930 -3885 970 -3875
rect 995 -3595 1035 -3585
rect 1810 -3510 1995 -3500
rect 1810 -3530 1890 -3510
rect 1910 -3530 1995 -3510
rect 1810 -3540 1995 -3530
rect 995 -3675 1000 -3595
rect 1020 -3675 1030 -3595
rect 995 -3795 1030 -3675
rect 995 -3875 1005 -3795
rect 1025 -3875 1030 -3795
rect 1810 -3695 1865 -3540
rect 2345 -3625 2375 -3380
rect 2458 -3415 2508 -3400
rect 2458 -3440 2473 -3415
rect 2493 -3440 2508 -3415
rect 2458 -3450 2508 -3440
rect 3435 -3485 3670 -3475
rect 2460 -3500 2500 -3490
rect 2460 -3580 2470 -3500
rect 2490 -3580 2500 -3500
rect 2460 -3625 2500 -3580
rect 1810 -3765 1820 -3695
rect 1850 -3765 1865 -3695
rect 1810 -3815 1865 -3765
rect 1925 -3695 1980 -3640
rect 2345 -3650 2500 -3625
rect 1925 -3765 1940 -3695
rect 1970 -3765 1980 -3695
rect 995 -3885 1030 -3875
rect 290 -3900 470 -3895
rect 135 -3920 175 -3915
rect 1815 -4020 1890 -4010
rect 1815 -4045 1840 -4020
rect 1870 -4045 1890 -4020
rect 1815 -4050 1890 -4045
rect 1925 -4065 1980 -3765
rect 2460 -3700 2500 -3650
rect 2460 -3780 2470 -3700
rect 2490 -3780 2500 -3700
rect 2460 -3790 2500 -3780
rect 2525 -3500 2560 -3490
rect 2525 -3580 2530 -3500
rect 2550 -3580 2560 -3500
rect 3435 -3510 3620 -3485
rect 3650 -3510 3670 -3485
rect 3435 -3515 3670 -3510
rect 2525 -3700 2560 -3580
rect 3705 -3530 3760 -3230
rect 4240 -3115 4250 -3095
rect 4270 -3115 4280 -3095
rect 4240 -3165 4280 -3115
rect 4240 -3245 4250 -3165
rect 4270 -3245 4280 -3165
rect 4240 -3255 4280 -3245
rect 4305 -2965 4340 -2955
rect 4305 -3045 4310 -2965
rect 4330 -3045 4340 -2965
rect 4305 -3165 4340 -3045
rect 4305 -3245 4315 -3165
rect 4335 -3245 4340 -3165
rect 6895 -2960 6975 -2940
rect 6995 -2960 7080 -2940
rect 6895 -2970 7080 -2960
rect 6895 -3125 6950 -2970
rect 7545 -3010 7555 -2930
rect 7575 -3010 7585 -2930
rect 7545 -3060 7585 -3010
rect 6895 -3195 6905 -3125
rect 6935 -3195 6950 -3125
rect 6895 -3245 6950 -3195
rect 7010 -3125 7065 -3070
rect 7010 -3195 7025 -3125
rect 7055 -3195 7065 -3125
rect 4305 -3340 4340 -3245
rect 4755 -3340 5680 -3315
rect 4305 -3345 5680 -3340
rect 4305 -3380 4775 -3345
rect 4233 -3475 4283 -3460
rect 4233 -3500 4248 -3475
rect 4268 -3500 4283 -3475
rect 4233 -3510 4283 -3500
rect 3980 -3525 4020 -3520
rect 3980 -3530 3990 -3525
rect 3705 -3550 3990 -3530
rect 4010 -3550 4020 -3525
rect 4305 -3550 4340 -3380
rect 4945 -3405 4995 -3390
rect 4945 -3430 4960 -3405
rect 4980 -3430 4995 -3405
rect 4945 -3440 4995 -3430
rect 2525 -3780 2535 -3700
rect 2555 -3780 2560 -3700
rect 2720 -3710 2770 -3695
rect 2720 -3735 2735 -3710
rect 2755 -3735 2770 -3710
rect 2720 -3745 2770 -3735
rect 3595 -3705 3645 -3695
rect 2525 -3875 2560 -3780
rect 2810 -3775 3015 -3765
rect 2810 -3800 2880 -3775
rect 2930 -3800 3015 -3775
rect 2810 -3810 3015 -3800
rect 3595 -3775 3605 -3705
rect 3635 -3775 3645 -3705
rect 2525 -3915 2755 -3875
rect 2453 -4010 2503 -3995
rect 2453 -4035 2468 -4010
rect 2488 -4035 2503 -4010
rect 2453 -4045 2503 -4035
rect 2200 -4060 2240 -4055
rect 2200 -4065 2210 -4060
rect 1925 -4085 2210 -4065
rect 2230 -4085 2240 -4060
rect 2525 -4085 2560 -3915
rect 883 -4175 933 -4160
rect 65 -4200 115 -4185
rect 65 -4225 80 -4200
rect 100 -4225 115 -4200
rect 883 -4200 898 -4175
rect 918 -4200 933 -4175
rect 883 -4210 933 -4200
rect 65 -4235 115 -4225
rect 1815 -4240 1865 -4230
rect 885 -4260 925 -4250
rect 235 -4270 420 -4260
rect 235 -4290 315 -4270
rect 335 -4290 420 -4270
rect 235 -4300 420 -4290
rect 235 -4455 290 -4300
rect 885 -4340 895 -4260
rect 915 -4340 925 -4260
rect 885 -4390 925 -4340
rect 235 -4525 245 -4455
rect 275 -4525 290 -4455
rect 235 -4575 290 -4525
rect 350 -4455 405 -4400
rect 350 -4525 365 -4455
rect 395 -4525 405 -4455
rect 95 -4780 315 -4770
rect 95 -4805 265 -4780
rect 295 -4805 315 -4780
rect 95 -4810 315 -4805
rect 350 -4825 405 -4525
rect 885 -4410 895 -4390
rect 915 -4410 925 -4390
rect 885 -4460 925 -4410
rect 885 -4540 895 -4460
rect 915 -4540 925 -4460
rect 885 -4550 925 -4540
rect 950 -4260 985 -4250
rect 950 -4340 955 -4260
rect 975 -4340 985 -4260
rect 950 -4460 985 -4340
rect 1815 -4310 1825 -4240
rect 1855 -4310 1865 -4240
rect 1815 -4350 1865 -4310
rect 1925 -4240 1980 -4085
rect 2200 -4090 2240 -4085
rect 2455 -4095 2495 -4085
rect 2455 -4175 2465 -4095
rect 2485 -4175 2495 -4095
rect 2455 -4230 2495 -4175
rect 1925 -4310 1935 -4240
rect 1965 -4310 1980 -4240
rect 1925 -4320 1980 -4310
rect 2240 -4260 2495 -4230
rect 1660 -4365 1865 -4350
rect 1660 -4375 1995 -4365
rect 1660 -4385 1885 -4375
rect 1660 -4390 1700 -4385
rect 1660 -4415 1670 -4390
rect 1690 -4415 1700 -4390
rect 1815 -4395 1885 -4385
rect 1910 -4395 1995 -4375
rect 1815 -4400 1995 -4395
rect 1660 -4420 1700 -4415
rect 950 -4540 960 -4460
rect 980 -4540 985 -4460
rect 950 -4630 985 -4540
rect 2240 -4630 2270 -4260
rect 2455 -4295 2495 -4260
rect 2455 -4375 2465 -4295
rect 2485 -4375 2495 -4295
rect 2455 -4385 2495 -4375
rect 2520 -4095 2560 -4085
rect 2520 -4175 2525 -4095
rect 2545 -4175 2555 -4095
rect 2520 -4295 2555 -4175
rect 2520 -4375 2530 -4295
rect 2550 -4375 2555 -4295
rect 2520 -4385 2555 -4375
rect 2725 -4385 2755 -3915
rect 2810 -3945 2890 -3810
rect 3595 -3815 3645 -3775
rect 3705 -3705 3760 -3550
rect 3980 -3555 4020 -3550
rect 3705 -3775 3715 -3705
rect 3745 -3775 3760 -3705
rect 3705 -3785 3760 -3775
rect 4235 -3560 4275 -3550
rect 4235 -3640 4245 -3560
rect 4265 -3640 4275 -3560
rect 4235 -3710 4275 -3640
rect 4235 -3730 4245 -3710
rect 4265 -3730 4275 -3710
rect 4235 -3760 4275 -3730
rect 3440 -3830 3645 -3815
rect 3440 -3840 3775 -3830
rect 3440 -3850 3665 -3840
rect 3440 -3855 3480 -3850
rect 3440 -3880 3450 -3855
rect 3470 -3880 3480 -3855
rect 3595 -3860 3665 -3850
rect 3690 -3860 3775 -3840
rect 4235 -3840 4245 -3760
rect 4265 -3840 4275 -3760
rect 4235 -3850 4275 -3840
rect 4300 -3560 4340 -3550
rect 5115 -3475 5300 -3465
rect 5115 -3495 5195 -3475
rect 5215 -3495 5300 -3475
rect 5115 -3505 5300 -3495
rect 4300 -3640 4305 -3560
rect 4325 -3640 4335 -3560
rect 4300 -3760 4335 -3640
rect 4300 -3840 4310 -3760
rect 4330 -3840 4335 -3760
rect 5115 -3660 5170 -3505
rect 5650 -3590 5680 -3345
rect 5763 -3380 5813 -3365
rect 5763 -3405 5778 -3380
rect 5798 -3405 5813 -3380
rect 5763 -3415 5813 -3405
rect 6740 -3450 6975 -3440
rect 5765 -3465 5805 -3455
rect 5765 -3545 5775 -3465
rect 5795 -3545 5805 -3465
rect 5765 -3590 5805 -3545
rect 5115 -3730 5125 -3660
rect 5155 -3730 5170 -3660
rect 5115 -3780 5170 -3730
rect 5230 -3660 5285 -3605
rect 5650 -3615 5805 -3590
rect 5230 -3730 5245 -3660
rect 5275 -3730 5285 -3660
rect 4300 -3850 4335 -3840
rect 3595 -3865 3775 -3860
rect 3440 -3885 3480 -3880
rect 2810 -4290 2820 -3945
rect 2885 -4290 2890 -3945
rect 2810 -4315 2890 -4290
rect 2930 -3945 3010 -3915
rect 2930 -4290 2935 -3945
rect 3000 -4290 3010 -3945
rect 5120 -3985 5195 -3975
rect 5120 -4010 5145 -3985
rect 5175 -4010 5195 -3985
rect 5120 -4015 5195 -4010
rect 5230 -4030 5285 -3730
rect 5765 -3665 5805 -3615
rect 5765 -3745 5775 -3665
rect 5795 -3745 5805 -3665
rect 5765 -3755 5805 -3745
rect 5830 -3465 5865 -3455
rect 5830 -3545 5835 -3465
rect 5855 -3545 5865 -3465
rect 6740 -3475 6925 -3450
rect 6955 -3475 6975 -3450
rect 6740 -3480 6975 -3475
rect 5830 -3665 5865 -3545
rect 7010 -3495 7065 -3195
rect 7545 -3080 7555 -3060
rect 7575 -3080 7585 -3060
rect 7545 -3130 7585 -3080
rect 7545 -3210 7555 -3130
rect 7575 -3210 7585 -3130
rect 7545 -3220 7585 -3210
rect 7610 -2930 7645 -2920
rect 7610 -3010 7615 -2930
rect 7635 -3010 7645 -2930
rect 7610 -3130 7645 -3010
rect 7610 -3210 7620 -3130
rect 7640 -3210 7645 -3130
rect 10200 -2925 10280 -2905
rect 10300 -2925 10385 -2905
rect 10200 -2935 10385 -2925
rect 10200 -3090 10255 -2935
rect 10850 -2975 10860 -2895
rect 10880 -2975 10890 -2895
rect 10850 -3025 10890 -2975
rect 10200 -3160 10210 -3090
rect 10240 -3160 10255 -3090
rect 10200 -3210 10255 -3160
rect 10315 -3090 10370 -3035
rect 10315 -3160 10330 -3090
rect 10360 -3160 10370 -3090
rect 7610 -3305 7645 -3210
rect 8060 -3305 8985 -3280
rect 7610 -3310 8985 -3305
rect 7610 -3345 8080 -3310
rect 7538 -3440 7588 -3425
rect 7538 -3465 7553 -3440
rect 7573 -3465 7588 -3440
rect 7538 -3475 7588 -3465
rect 7285 -3490 7325 -3485
rect 7285 -3495 7295 -3490
rect 7010 -3515 7295 -3495
rect 7315 -3515 7325 -3490
rect 7610 -3515 7645 -3345
rect 8250 -3370 8300 -3355
rect 8250 -3395 8265 -3370
rect 8285 -3395 8300 -3370
rect 8250 -3405 8300 -3395
rect 5830 -3745 5840 -3665
rect 5860 -3745 5865 -3665
rect 6050 -3675 6100 -3660
rect 6050 -3700 6065 -3675
rect 6085 -3700 6100 -3675
rect 6050 -3710 6100 -3700
rect 6900 -3670 6950 -3660
rect 5830 -3840 5865 -3745
rect 6140 -3740 6345 -3730
rect 6140 -3765 6210 -3740
rect 6260 -3765 6345 -3740
rect 6140 -3775 6345 -3765
rect 6900 -3740 6910 -3670
rect 6940 -3740 6950 -3670
rect 5830 -3880 6085 -3840
rect 5758 -3975 5808 -3960
rect 5758 -4000 5773 -3975
rect 5793 -4000 5808 -3975
rect 5758 -4010 5808 -4000
rect 5505 -4025 5545 -4020
rect 5505 -4030 5515 -4025
rect 5230 -4050 5515 -4030
rect 5535 -4050 5545 -4025
rect 5830 -4050 5865 -3880
rect 4188 -4140 4238 -4125
rect 3370 -4165 3420 -4150
rect 3370 -4190 3385 -4165
rect 3405 -4190 3420 -4165
rect 4188 -4165 4203 -4140
rect 4223 -4165 4238 -4140
rect 4188 -4175 4238 -4165
rect 3370 -4200 3420 -4190
rect 5120 -4205 5170 -4195
rect 4190 -4225 4230 -4215
rect 2930 -4365 3010 -4290
rect 3540 -4235 3725 -4225
rect 3540 -4255 3620 -4235
rect 3640 -4255 3725 -4235
rect 3540 -4265 3725 -4255
rect 2725 -4395 2900 -4385
rect 2725 -4415 2870 -4395
rect 2890 -4415 2900 -4395
rect 2725 -4425 2900 -4415
rect 2930 -4425 3115 -4365
rect 950 -4675 2270 -4630
rect 2810 -4545 2890 -4515
rect 878 -4770 928 -4755
rect 878 -4795 893 -4770
rect 913 -4795 928 -4770
rect 878 -4805 928 -4795
rect 625 -4820 665 -4815
rect 625 -4825 635 -4820
rect 350 -4845 635 -4825
rect 655 -4845 665 -4820
rect 950 -4845 985 -4675
rect 2810 -4700 2820 -4545
rect 2875 -4700 2890 -4545
rect 2655 -4730 2890 -4700
rect 2930 -4545 3010 -4425
rect 2930 -4700 2945 -4545
rect 3000 -4700 3010 -4545
rect 2930 -4715 3010 -4700
rect 2655 -4735 2750 -4730
rect 2655 -4740 2695 -4735
rect 2655 -4765 2665 -4740
rect 2685 -4765 2695 -4740
rect 2655 -4770 2695 -4765
rect 2810 -4755 2890 -4730
rect 2810 -4775 2825 -4755
rect 2865 -4775 2890 -4755
rect 2810 -4785 2890 -4775
rect 240 -5000 290 -4990
rect 240 -5070 250 -5000
rect 280 -5070 290 -5000
rect 240 -5110 290 -5070
rect 350 -5000 405 -4845
rect 625 -4850 665 -4845
rect 350 -5070 360 -5000
rect 390 -5070 405 -5000
rect 350 -5080 405 -5070
rect 880 -4855 920 -4845
rect 880 -4935 890 -4855
rect 910 -4935 920 -4855
rect 880 -5005 920 -4935
rect 880 -5025 890 -5005
rect 910 -5025 920 -5005
rect 880 -5055 920 -5025
rect 85 -5125 290 -5110
rect 85 -5135 420 -5125
rect 85 -5145 310 -5135
rect 85 -5150 125 -5145
rect 85 -5175 95 -5150
rect 115 -5175 125 -5150
rect 240 -5155 310 -5145
rect 335 -5155 420 -5135
rect 880 -5135 890 -5055
rect 910 -5135 920 -5055
rect 880 -5145 920 -5135
rect 945 -4855 985 -4845
rect 945 -4935 950 -4855
rect 970 -4935 980 -4855
rect 3065 -4915 3115 -4425
rect 3540 -4420 3595 -4265
rect 4190 -4305 4200 -4225
rect 4220 -4305 4230 -4225
rect 4190 -4355 4230 -4305
rect 3540 -4490 3550 -4420
rect 3580 -4490 3595 -4420
rect 3540 -4540 3595 -4490
rect 3655 -4420 3710 -4365
rect 3655 -4490 3670 -4420
rect 3700 -4490 3710 -4420
rect 3400 -4745 3620 -4735
rect 3400 -4770 3570 -4745
rect 3600 -4770 3620 -4745
rect 3400 -4775 3620 -4770
rect 945 -5055 980 -4935
rect 945 -5135 955 -5055
rect 975 -5135 980 -5055
rect 945 -5145 980 -5135
rect 2670 -4965 3115 -4915
rect 3655 -4790 3710 -4490
rect 4190 -4375 4200 -4355
rect 4220 -4375 4230 -4355
rect 4190 -4425 4230 -4375
rect 4190 -4505 4200 -4425
rect 4220 -4505 4230 -4425
rect 4190 -4515 4230 -4505
rect 4255 -4225 4290 -4215
rect 4255 -4305 4260 -4225
rect 4280 -4305 4290 -4225
rect 4255 -4425 4290 -4305
rect 5120 -4275 5130 -4205
rect 5160 -4275 5170 -4205
rect 5120 -4315 5170 -4275
rect 5230 -4205 5285 -4050
rect 5505 -4055 5545 -4050
rect 5760 -4060 5800 -4050
rect 5760 -4140 5770 -4060
rect 5790 -4140 5800 -4060
rect 5760 -4195 5800 -4140
rect 5230 -4275 5240 -4205
rect 5270 -4275 5285 -4205
rect 5230 -4285 5285 -4275
rect 5545 -4225 5800 -4195
rect 4965 -4330 5170 -4315
rect 4965 -4340 5300 -4330
rect 4965 -4350 5190 -4340
rect 4965 -4355 5005 -4350
rect 4965 -4380 4975 -4355
rect 4995 -4380 5005 -4355
rect 5120 -4360 5190 -4350
rect 5215 -4360 5300 -4340
rect 5120 -4365 5300 -4360
rect 4965 -4385 5005 -4380
rect 4255 -4505 4265 -4425
rect 4285 -4505 4290 -4425
rect 4255 -4590 4290 -4505
rect 4255 -4595 4460 -4590
rect 5545 -4595 5575 -4225
rect 5760 -4260 5800 -4225
rect 5760 -4340 5770 -4260
rect 5790 -4340 5800 -4260
rect 5760 -4350 5800 -4340
rect 5825 -4060 5865 -4050
rect 5825 -4140 5830 -4060
rect 5850 -4140 5860 -4060
rect 5825 -4260 5860 -4140
rect 5825 -4340 5835 -4260
rect 5855 -4340 5860 -4260
rect 5825 -4350 5860 -4340
rect 6055 -4350 6085 -3880
rect 6140 -3910 6220 -3775
rect 6900 -3780 6950 -3740
rect 7010 -3670 7065 -3515
rect 7285 -3520 7325 -3515
rect 7010 -3740 7020 -3670
rect 7050 -3740 7065 -3670
rect 7010 -3750 7065 -3740
rect 7540 -3525 7580 -3515
rect 7540 -3605 7550 -3525
rect 7570 -3605 7580 -3525
rect 7540 -3675 7580 -3605
rect 7540 -3695 7550 -3675
rect 7570 -3695 7580 -3675
rect 7540 -3725 7580 -3695
rect 6745 -3795 6950 -3780
rect 6745 -3805 7080 -3795
rect 6745 -3815 6970 -3805
rect 6745 -3820 6785 -3815
rect 6745 -3845 6755 -3820
rect 6775 -3845 6785 -3820
rect 6900 -3825 6970 -3815
rect 6995 -3825 7080 -3805
rect 7540 -3805 7550 -3725
rect 7570 -3805 7580 -3725
rect 7540 -3815 7580 -3805
rect 7605 -3525 7645 -3515
rect 8420 -3440 8605 -3430
rect 8420 -3460 8500 -3440
rect 8520 -3460 8605 -3440
rect 8420 -3470 8605 -3460
rect 7605 -3605 7610 -3525
rect 7630 -3605 7640 -3525
rect 7605 -3725 7640 -3605
rect 7605 -3805 7615 -3725
rect 7635 -3805 7640 -3725
rect 8420 -3625 8475 -3470
rect 8955 -3555 8985 -3310
rect 9068 -3345 9118 -3330
rect 9068 -3370 9083 -3345
rect 9103 -3370 9118 -3345
rect 9068 -3380 9118 -3370
rect 10045 -3415 10280 -3405
rect 9070 -3430 9110 -3420
rect 9070 -3510 9080 -3430
rect 9100 -3510 9110 -3430
rect 9070 -3555 9110 -3510
rect 8420 -3695 8430 -3625
rect 8460 -3695 8475 -3625
rect 8420 -3745 8475 -3695
rect 8535 -3625 8590 -3570
rect 8955 -3580 9110 -3555
rect 8535 -3695 8550 -3625
rect 8580 -3695 8590 -3625
rect 7605 -3815 7640 -3805
rect 6900 -3830 7080 -3825
rect 6745 -3850 6785 -3845
rect 6140 -4255 6150 -3910
rect 6215 -4255 6220 -3910
rect 6140 -4280 6220 -4255
rect 6260 -3910 6340 -3880
rect 6260 -4255 6265 -3910
rect 6330 -4255 6340 -3910
rect 8425 -3950 8500 -3940
rect 8425 -3975 8450 -3950
rect 8480 -3975 8500 -3950
rect 8425 -3980 8500 -3975
rect 8535 -3995 8590 -3695
rect 9070 -3630 9110 -3580
rect 9070 -3710 9080 -3630
rect 9100 -3710 9110 -3630
rect 9070 -3720 9110 -3710
rect 9135 -3430 9170 -3420
rect 9135 -3510 9140 -3430
rect 9160 -3510 9170 -3430
rect 10045 -3440 10230 -3415
rect 10260 -3440 10280 -3415
rect 10045 -3445 10280 -3440
rect 9135 -3630 9170 -3510
rect 10315 -3460 10370 -3160
rect 10850 -3045 10860 -3025
rect 10880 -3045 10890 -3025
rect 10850 -3095 10890 -3045
rect 10850 -3175 10860 -3095
rect 10880 -3175 10890 -3095
rect 10850 -3185 10890 -3175
rect 10915 -2895 10950 -2885
rect 10915 -2975 10920 -2895
rect 10940 -2975 10950 -2895
rect 10915 -3095 10950 -2975
rect 13635 -3065 13685 -3050
rect 13635 -3090 13650 -3065
rect 13670 -3090 13685 -3065
rect 10915 -3175 10925 -3095
rect 10945 -3175 10950 -3095
rect 13205 -3105 13255 -3090
rect 13635 -3100 13685 -3090
rect 13205 -3130 13220 -3105
rect 13240 -3130 13255 -3105
rect 13205 -3140 13255 -3130
rect 13725 -3130 13930 -3120
rect 13725 -3155 13795 -3130
rect 13845 -3155 13930 -3130
rect 10915 -3270 10950 -3175
rect 13295 -3170 13500 -3160
rect 13295 -3195 13365 -3170
rect 13415 -3195 13500 -3170
rect 13295 -3205 13500 -3195
rect 13725 -3165 13930 -3155
rect 11365 -3270 12290 -3245
rect 10915 -3275 12290 -3270
rect 10915 -3310 11385 -3275
rect 10843 -3405 10893 -3390
rect 10843 -3430 10858 -3405
rect 10878 -3430 10893 -3405
rect 10843 -3440 10893 -3430
rect 10590 -3455 10630 -3450
rect 10590 -3460 10600 -3455
rect 10315 -3480 10600 -3460
rect 10620 -3480 10630 -3455
rect 10915 -3480 10950 -3310
rect 11555 -3335 11605 -3320
rect 11555 -3360 11570 -3335
rect 11590 -3360 11605 -3335
rect 11555 -3370 11605 -3360
rect 9135 -3710 9145 -3630
rect 9165 -3710 9170 -3630
rect 9365 -3640 9415 -3625
rect 9365 -3665 9380 -3640
rect 9400 -3665 9415 -3640
rect 9365 -3675 9415 -3665
rect 10205 -3635 10255 -3625
rect 9135 -3805 9170 -3710
rect 9455 -3705 9660 -3695
rect 9455 -3730 9525 -3705
rect 9575 -3730 9660 -3705
rect 9455 -3740 9660 -3730
rect 10205 -3705 10215 -3635
rect 10245 -3705 10255 -3635
rect 9135 -3845 9400 -3805
rect 9063 -3940 9113 -3925
rect 9063 -3965 9078 -3940
rect 9098 -3965 9113 -3940
rect 9063 -3975 9113 -3965
rect 8810 -3990 8850 -3985
rect 8810 -3995 8820 -3990
rect 8535 -4015 8820 -3995
rect 8840 -4015 8850 -3990
rect 9135 -4015 9170 -3845
rect 7493 -4105 7543 -4090
rect 6675 -4130 6725 -4115
rect 6675 -4155 6690 -4130
rect 6710 -4155 6725 -4130
rect 7493 -4130 7508 -4105
rect 7528 -4130 7543 -4105
rect 7493 -4140 7543 -4130
rect 6675 -4165 6725 -4155
rect 8425 -4170 8475 -4160
rect 7495 -4190 7535 -4180
rect 6260 -4345 6340 -4255
rect 6845 -4200 7030 -4190
rect 6845 -4220 6925 -4200
rect 6945 -4220 7030 -4200
rect 6845 -4230 7030 -4220
rect 6055 -4360 6230 -4350
rect 6055 -4380 6200 -4360
rect 6220 -4380 6230 -4360
rect 6055 -4390 6230 -4380
rect 6260 -4405 6450 -4345
rect 4255 -4640 5575 -4595
rect 6140 -4510 6220 -4480
rect 4183 -4735 4233 -4720
rect 4183 -4760 4198 -4735
rect 4218 -4760 4233 -4735
rect 4183 -4770 4233 -4760
rect 3930 -4785 3970 -4780
rect 3930 -4790 3940 -4785
rect 3655 -4810 3940 -4790
rect 3960 -4810 3970 -4785
rect 4255 -4810 4290 -4640
rect 6140 -4665 6150 -4510
rect 6205 -4665 6220 -4510
rect 5985 -4695 6220 -4665
rect 6260 -4510 6340 -4405
rect 6260 -4665 6275 -4510
rect 6330 -4665 6340 -4510
rect 6260 -4680 6340 -4665
rect 5985 -4700 6080 -4695
rect 5985 -4705 6025 -4700
rect 5985 -4730 5995 -4705
rect 6015 -4730 6025 -4705
rect 5985 -4735 6025 -4730
rect 6140 -4720 6220 -4695
rect 6140 -4740 6155 -4720
rect 6195 -4740 6220 -4720
rect 6140 -4750 6220 -4740
rect 3545 -4965 3595 -4955
rect 240 -5160 420 -5155
rect 85 -5180 125 -5175
rect 2670 -5695 2715 -4965
rect 3545 -5035 3555 -4965
rect 3585 -5035 3595 -4965
rect 3545 -5075 3595 -5035
rect 3655 -4965 3710 -4810
rect 3930 -4815 3970 -4810
rect 3655 -5035 3665 -4965
rect 3695 -5035 3710 -4965
rect 3655 -5045 3710 -5035
rect 4185 -4820 4225 -4810
rect 4185 -4900 4195 -4820
rect 4215 -4900 4225 -4820
rect 4185 -4970 4225 -4900
rect 4185 -4990 4195 -4970
rect 4215 -4990 4225 -4970
rect 4185 -5020 4225 -4990
rect 3390 -5090 3595 -5075
rect 3390 -5100 3725 -5090
rect 3390 -5110 3615 -5100
rect 3390 -5115 3430 -5110
rect 3390 -5140 3400 -5115
rect 3420 -5140 3430 -5115
rect 3545 -5120 3615 -5110
rect 3640 -5120 3725 -5100
rect 4185 -5100 4195 -5020
rect 4215 -5100 4225 -5020
rect 4185 -5110 4225 -5100
rect 4250 -4820 4290 -4810
rect 4250 -4900 4255 -4820
rect 4275 -4900 4285 -4820
rect 6415 -4895 6450 -4405
rect 6845 -4385 6900 -4230
rect 7495 -4270 7505 -4190
rect 7525 -4270 7535 -4190
rect 7495 -4320 7535 -4270
rect 6845 -4455 6855 -4385
rect 6885 -4455 6900 -4385
rect 6845 -4505 6900 -4455
rect 6960 -4385 7015 -4330
rect 6960 -4455 6975 -4385
rect 7005 -4455 7015 -4385
rect 6705 -4710 6925 -4700
rect 6705 -4735 6875 -4710
rect 6905 -4735 6925 -4710
rect 6705 -4740 6925 -4735
rect 4250 -5020 4285 -4900
rect 4250 -5100 4260 -5020
rect 4280 -5100 4285 -5020
rect 4250 -5110 4285 -5100
rect 6125 -4950 6450 -4895
rect 6960 -4755 7015 -4455
rect 7495 -4340 7505 -4320
rect 7525 -4340 7535 -4320
rect 7495 -4390 7535 -4340
rect 7495 -4470 7505 -4390
rect 7525 -4470 7535 -4390
rect 7495 -4480 7535 -4470
rect 7560 -4190 7595 -4180
rect 7560 -4270 7565 -4190
rect 7585 -4270 7595 -4190
rect 7560 -4390 7595 -4270
rect 8425 -4240 8435 -4170
rect 8465 -4240 8475 -4170
rect 8425 -4280 8475 -4240
rect 8535 -4170 8590 -4015
rect 8810 -4020 8850 -4015
rect 9065 -4025 9105 -4015
rect 9065 -4105 9075 -4025
rect 9095 -4105 9105 -4025
rect 9065 -4160 9105 -4105
rect 8535 -4240 8545 -4170
rect 8575 -4240 8590 -4170
rect 8535 -4250 8590 -4240
rect 8850 -4190 9105 -4160
rect 8270 -4295 8475 -4280
rect 8270 -4305 8605 -4295
rect 8270 -4315 8495 -4305
rect 8270 -4320 8310 -4315
rect 8270 -4345 8280 -4320
rect 8300 -4345 8310 -4320
rect 8425 -4325 8495 -4315
rect 8520 -4325 8605 -4305
rect 8425 -4330 8605 -4325
rect 8270 -4350 8310 -4345
rect 7560 -4470 7570 -4390
rect 7590 -4470 7595 -4390
rect 7560 -4555 7595 -4470
rect 7560 -4560 7765 -4555
rect 8850 -4560 8880 -4190
rect 9065 -4225 9105 -4190
rect 9065 -4305 9075 -4225
rect 9095 -4305 9105 -4225
rect 9065 -4315 9105 -4305
rect 9130 -4025 9170 -4015
rect 9130 -4105 9135 -4025
rect 9155 -4105 9165 -4025
rect 9130 -4225 9165 -4105
rect 9130 -4305 9140 -4225
rect 9160 -4305 9165 -4225
rect 9130 -4315 9165 -4305
rect 9370 -4315 9400 -3845
rect 9455 -3875 9535 -3740
rect 10205 -3745 10255 -3705
rect 10315 -3635 10370 -3480
rect 10590 -3485 10630 -3480
rect 10315 -3705 10325 -3635
rect 10355 -3705 10370 -3635
rect 10315 -3715 10370 -3705
rect 10845 -3490 10885 -3480
rect 10845 -3570 10855 -3490
rect 10875 -3570 10885 -3490
rect 10845 -3640 10885 -3570
rect 10845 -3660 10855 -3640
rect 10875 -3660 10885 -3640
rect 10845 -3690 10885 -3660
rect 10050 -3760 10255 -3745
rect 10050 -3770 10385 -3760
rect 10050 -3780 10275 -3770
rect 10050 -3785 10090 -3780
rect 10050 -3810 10060 -3785
rect 10080 -3810 10090 -3785
rect 10205 -3790 10275 -3780
rect 10300 -3790 10385 -3770
rect 10845 -3770 10855 -3690
rect 10875 -3770 10885 -3690
rect 10845 -3780 10885 -3770
rect 10910 -3490 10950 -3480
rect 11725 -3405 11910 -3395
rect 11725 -3425 11805 -3405
rect 11825 -3425 11910 -3405
rect 11725 -3435 11910 -3425
rect 10910 -3570 10915 -3490
rect 10935 -3570 10945 -3490
rect 10910 -3690 10945 -3570
rect 10910 -3770 10920 -3690
rect 10940 -3770 10945 -3690
rect 11725 -3590 11780 -3435
rect 12260 -3520 12290 -3275
rect 12373 -3310 12423 -3295
rect 12373 -3335 12388 -3310
rect 12408 -3335 12423 -3310
rect 12373 -3345 12423 -3335
rect 13295 -3340 13375 -3205
rect 13725 -3300 13805 -3165
rect 12375 -3395 12415 -3385
rect 12375 -3475 12385 -3395
rect 12405 -3475 12415 -3395
rect 12375 -3520 12415 -3475
rect 11725 -3660 11735 -3590
rect 11765 -3660 11780 -3590
rect 11725 -3710 11780 -3660
rect 11840 -3590 11895 -3535
rect 12260 -3545 12415 -3520
rect 11840 -3660 11855 -3590
rect 11885 -3660 11895 -3590
rect 10910 -3780 10945 -3770
rect 10205 -3795 10385 -3790
rect 10050 -3815 10090 -3810
rect 9455 -4220 9465 -3875
rect 9530 -4220 9535 -3875
rect 9455 -4245 9535 -4220
rect 9575 -3875 9655 -3845
rect 9575 -4220 9580 -3875
rect 9645 -4220 9655 -3875
rect 11730 -3915 11805 -3905
rect 11730 -3940 11755 -3915
rect 11785 -3940 11805 -3915
rect 11730 -3945 11805 -3940
rect 11840 -3960 11895 -3660
rect 12375 -3595 12415 -3545
rect 12375 -3675 12385 -3595
rect 12405 -3675 12415 -3595
rect 12375 -3685 12415 -3675
rect 12440 -3395 12475 -3385
rect 12440 -3475 12445 -3395
rect 12465 -3475 12475 -3395
rect 12440 -3595 12475 -3475
rect 12440 -3675 12450 -3595
rect 12470 -3675 12475 -3595
rect 12440 -3770 12475 -3675
rect 13295 -3685 13305 -3340
rect 13370 -3685 13375 -3340
rect 13295 -3710 13375 -3685
rect 13415 -3340 13495 -3310
rect 13415 -3685 13420 -3340
rect 13485 -3685 13495 -3340
rect 13725 -3645 13735 -3300
rect 13800 -3645 13805 -3300
rect 13725 -3670 13805 -3645
rect 13845 -3300 13925 -3270
rect 13845 -3645 13850 -3300
rect 13915 -3645 13925 -3300
rect 13415 -3740 13495 -3685
rect 13415 -3750 13815 -3740
rect 13415 -3770 13785 -3750
rect 13805 -3770 13815 -3750
rect 12440 -3780 13255 -3770
rect 13415 -3780 13815 -3770
rect 12440 -3790 13385 -3780
rect 12440 -3810 13355 -3790
rect 13375 -3810 13385 -3790
rect 12368 -3905 12418 -3890
rect 12368 -3930 12383 -3905
rect 12403 -3930 12418 -3905
rect 12368 -3940 12418 -3930
rect 12115 -3955 12155 -3950
rect 12115 -3960 12125 -3955
rect 11840 -3980 12125 -3960
rect 12145 -3980 12155 -3955
rect 12440 -3980 12475 -3810
rect 13240 -3820 13385 -3810
rect 10798 -4070 10848 -4055
rect 9980 -4095 10030 -4080
rect 9980 -4120 9995 -4095
rect 10015 -4120 10030 -4095
rect 10798 -4095 10813 -4070
rect 10833 -4095 10848 -4070
rect 10798 -4105 10848 -4095
rect 9980 -4130 10030 -4120
rect 11730 -4135 11780 -4125
rect 10800 -4155 10840 -4145
rect 9575 -4315 9655 -4220
rect 10150 -4165 10335 -4155
rect 10150 -4185 10230 -4165
rect 10250 -4185 10335 -4165
rect 10150 -4195 10335 -4185
rect 9370 -4325 9545 -4315
rect 9370 -4345 9515 -4325
rect 9535 -4345 9545 -4325
rect 9370 -4355 9545 -4345
rect 9575 -4375 9740 -4315
rect 7560 -4605 8880 -4560
rect 9455 -4475 9535 -4445
rect 7488 -4700 7538 -4685
rect 7488 -4725 7503 -4700
rect 7523 -4725 7538 -4700
rect 7488 -4735 7538 -4725
rect 7235 -4750 7275 -4745
rect 7235 -4755 7245 -4750
rect 6960 -4775 7245 -4755
rect 7265 -4775 7275 -4750
rect 7560 -4775 7595 -4605
rect 9455 -4630 9465 -4475
rect 9520 -4630 9535 -4475
rect 9300 -4660 9535 -4630
rect 9575 -4475 9655 -4375
rect 9575 -4630 9590 -4475
rect 9645 -4630 9655 -4475
rect 9575 -4645 9655 -4630
rect 9300 -4665 9395 -4660
rect 9300 -4670 9340 -4665
rect 9300 -4695 9310 -4670
rect 9330 -4695 9340 -4670
rect 9300 -4700 9340 -4695
rect 9455 -4685 9535 -4660
rect 9455 -4705 9470 -4685
rect 9510 -4705 9535 -4685
rect 9455 -4715 9535 -4705
rect 6850 -4930 6900 -4920
rect 3545 -5125 3725 -5120
rect 3390 -5145 3430 -5140
rect 2795 -5530 2845 -5515
rect 2795 -5555 2810 -5530
rect 2830 -5555 2845 -5530
rect 2795 -5565 2845 -5555
rect 2885 -5595 3090 -5585
rect 2885 -5620 2955 -5595
rect 3005 -5620 3090 -5595
rect 2885 -5630 3090 -5620
rect 6125 -5590 6180 -4950
rect 6850 -5000 6860 -4930
rect 6890 -5000 6900 -4930
rect 6850 -5040 6900 -5000
rect 6960 -4930 7015 -4775
rect 7235 -4780 7275 -4775
rect 6960 -5000 6970 -4930
rect 7000 -5000 7015 -4930
rect 6960 -5010 7015 -5000
rect 7490 -4785 7530 -4775
rect 7490 -4865 7500 -4785
rect 7520 -4865 7530 -4785
rect 7490 -4935 7530 -4865
rect 7490 -4955 7500 -4935
rect 7520 -4955 7530 -4935
rect 7490 -4985 7530 -4955
rect 6695 -5055 6900 -5040
rect 6695 -5065 7030 -5055
rect 6695 -5075 6920 -5065
rect 6695 -5080 6735 -5075
rect 6695 -5105 6705 -5080
rect 6725 -5105 6735 -5080
rect 6850 -5085 6920 -5075
rect 6945 -5085 7030 -5065
rect 7490 -5065 7500 -4985
rect 7520 -5065 7530 -4985
rect 7490 -5075 7530 -5065
rect 7555 -4785 7595 -4775
rect 7555 -4865 7560 -4785
rect 7580 -4865 7590 -4785
rect 7555 -4985 7590 -4865
rect 9700 -4870 9740 -4375
rect 10150 -4350 10205 -4195
rect 10800 -4235 10810 -4155
rect 10830 -4235 10840 -4155
rect 10800 -4285 10840 -4235
rect 10150 -4420 10160 -4350
rect 10190 -4420 10205 -4350
rect 10150 -4470 10205 -4420
rect 10265 -4350 10320 -4295
rect 10265 -4420 10280 -4350
rect 10310 -4420 10320 -4350
rect 10010 -4675 10230 -4665
rect 10010 -4700 10180 -4675
rect 10210 -4700 10230 -4675
rect 10010 -4705 10230 -4700
rect 7555 -5065 7565 -4985
rect 7585 -5065 7590 -4985
rect 7555 -5075 7590 -5065
rect 9230 -4915 9740 -4870
rect 10265 -4720 10320 -4420
rect 10800 -4305 10810 -4285
rect 10830 -4305 10840 -4285
rect 10800 -4355 10840 -4305
rect 10800 -4435 10810 -4355
rect 10830 -4435 10840 -4355
rect 10800 -4445 10840 -4435
rect 10865 -4155 10900 -4145
rect 10865 -4235 10870 -4155
rect 10890 -4235 10900 -4155
rect 10865 -4355 10900 -4235
rect 11730 -4205 11740 -4135
rect 11770 -4205 11780 -4135
rect 11730 -4245 11780 -4205
rect 11840 -4135 11895 -3980
rect 12115 -3985 12155 -3980
rect 12370 -3990 12410 -3980
rect 12370 -4070 12380 -3990
rect 12400 -4070 12410 -3990
rect 12370 -4125 12410 -4070
rect 11840 -4205 11850 -4135
rect 11880 -4205 11895 -4135
rect 11840 -4215 11895 -4205
rect 12155 -4155 12410 -4125
rect 11575 -4260 11780 -4245
rect 11575 -4270 11910 -4260
rect 11575 -4280 11800 -4270
rect 11575 -4285 11615 -4280
rect 11575 -4310 11585 -4285
rect 11605 -4310 11615 -4285
rect 11730 -4290 11800 -4280
rect 11825 -4290 11910 -4270
rect 11730 -4295 11910 -4290
rect 11575 -4315 11615 -4310
rect 10865 -4435 10875 -4355
rect 10895 -4435 10900 -4355
rect 10865 -4520 10900 -4435
rect 10865 -4525 11070 -4520
rect 12155 -4525 12185 -4155
rect 12370 -4190 12410 -4155
rect 12370 -4270 12380 -4190
rect 12400 -4270 12410 -4190
rect 12370 -4280 12410 -4270
rect 12435 -3990 12475 -3980
rect 13295 -3940 13375 -3910
rect 12435 -4070 12440 -3990
rect 12460 -4070 12470 -3990
rect 12435 -4190 12470 -4070
rect 13295 -4095 13305 -3940
rect 13360 -4095 13375 -3940
rect 13140 -4125 13375 -4095
rect 13415 -3940 13495 -3780
rect 13415 -4095 13430 -3940
rect 13485 -4095 13495 -3940
rect 13725 -3900 13805 -3870
rect 13725 -4055 13735 -3900
rect 13790 -4055 13805 -3900
rect 13415 -4110 13495 -4095
rect 13570 -4085 13805 -4055
rect 13845 -3900 13925 -3645
rect 13845 -4055 13860 -3900
rect 13915 -4055 13925 -3900
rect 13845 -4070 13925 -4055
rect 13570 -4090 13665 -4085
rect 13570 -4095 13610 -4090
rect 13570 -4120 13580 -4095
rect 13600 -4120 13610 -4095
rect 13570 -4125 13610 -4120
rect 13725 -4110 13805 -4085
rect 13140 -4130 13235 -4125
rect 13140 -4135 13180 -4130
rect 13140 -4160 13150 -4135
rect 13170 -4160 13180 -4135
rect 13140 -4165 13180 -4160
rect 13295 -4150 13375 -4125
rect 13725 -4130 13740 -4110
rect 13780 -4130 13805 -4110
rect 13725 -4140 13805 -4130
rect 13295 -4170 13310 -4150
rect 13350 -4170 13375 -4150
rect 13295 -4180 13375 -4170
rect 12435 -4270 12445 -4190
rect 12465 -4270 12470 -4190
rect 12435 -4280 12470 -4270
rect 10865 -4570 12185 -4525
rect 10793 -4665 10843 -4650
rect 10793 -4690 10808 -4665
rect 10828 -4690 10843 -4665
rect 10793 -4700 10843 -4690
rect 10540 -4715 10580 -4710
rect 10540 -4720 10550 -4715
rect 10265 -4740 10550 -4720
rect 10570 -4740 10580 -4715
rect 10865 -4740 10900 -4570
rect 10155 -4895 10205 -4885
rect 6850 -5090 7030 -5085
rect 6695 -5110 6735 -5105
rect 6240 -5425 6290 -5410
rect 6240 -5450 6255 -5425
rect 6275 -5450 6290 -5425
rect 6240 -5460 6290 -5450
rect 9230 -5470 9275 -4915
rect 10155 -4965 10165 -4895
rect 10195 -4965 10205 -4895
rect 10155 -5005 10205 -4965
rect 10265 -4895 10320 -4740
rect 10540 -4745 10580 -4740
rect 10265 -4965 10275 -4895
rect 10305 -4965 10320 -4895
rect 10265 -4975 10320 -4965
rect 10795 -4750 10835 -4740
rect 10795 -4830 10805 -4750
rect 10825 -4830 10835 -4750
rect 10795 -4900 10835 -4830
rect 10795 -4920 10805 -4900
rect 10825 -4920 10835 -4900
rect 10795 -4950 10835 -4920
rect 10000 -5020 10205 -5005
rect 10000 -5030 10335 -5020
rect 10000 -5040 10225 -5030
rect 10000 -5045 10040 -5040
rect 10000 -5070 10010 -5045
rect 10030 -5070 10040 -5045
rect 10155 -5050 10225 -5040
rect 10250 -5050 10335 -5030
rect 10795 -5030 10805 -4950
rect 10825 -5030 10835 -4950
rect 10795 -5040 10835 -5030
rect 10860 -4750 10900 -4740
rect 10860 -4830 10865 -4750
rect 10885 -4830 10895 -4750
rect 10860 -4950 10895 -4830
rect 10860 -5030 10870 -4950
rect 10890 -5030 10895 -4950
rect 10860 -5040 10895 -5030
rect 10155 -5055 10335 -5050
rect 10000 -5075 10040 -5070
rect 9345 -5305 9395 -5290
rect 9345 -5330 9360 -5305
rect 9380 -5330 9395 -5305
rect 9345 -5340 9395 -5330
rect 9435 -5370 9640 -5360
rect 9435 -5395 9505 -5370
rect 9555 -5395 9640 -5370
rect 9435 -5405 9640 -5395
rect 6330 -5490 6535 -5480
rect 6330 -5515 6400 -5490
rect 6450 -5515 6535 -5490
rect 9230 -5510 9380 -5470
rect 6330 -5525 6535 -5515
rect 6125 -5630 6275 -5590
rect 2670 -5735 2830 -5695
rect 2800 -6205 2830 -5735
rect 2885 -5765 2965 -5630
rect 2885 -6110 2895 -5765
rect 2960 -6110 2965 -5765
rect 2885 -6135 2965 -6110
rect 3005 -5765 3085 -5735
rect 3005 -6110 3010 -5765
rect 3075 -6110 3085 -5765
rect 2800 -6215 2975 -6205
rect 2800 -6235 2945 -6215
rect 2965 -6235 2975 -6215
rect 2800 -6245 2975 -6235
rect 2885 -6365 2965 -6335
rect 2885 -6520 2895 -6365
rect 2950 -6520 2965 -6365
rect 2730 -6550 2965 -6520
rect 3005 -6365 3085 -6110
rect 6245 -6100 6275 -5630
rect 6330 -5660 6410 -5525
rect 6330 -6005 6340 -5660
rect 6405 -6005 6410 -5660
rect 6330 -6030 6410 -6005
rect 6450 -5660 6530 -5630
rect 6450 -6005 6455 -5660
rect 6520 -6005 6530 -5660
rect 6245 -6110 6420 -6100
rect 6245 -6130 6390 -6110
rect 6410 -6130 6420 -6110
rect 6245 -6140 6420 -6130
rect 3005 -6520 3020 -6365
rect 3075 -6520 3085 -6365
rect 6330 -6260 6410 -6230
rect 6330 -6415 6340 -6260
rect 6395 -6415 6410 -6260
rect 6175 -6445 6410 -6415
rect 6450 -6260 6530 -6005
rect 9350 -5980 9380 -5510
rect 9435 -5540 9515 -5405
rect 9435 -5885 9445 -5540
rect 9510 -5885 9515 -5540
rect 9435 -5910 9515 -5885
rect 9555 -5540 9635 -5510
rect 9555 -5885 9560 -5540
rect 9625 -5885 9635 -5540
rect 9350 -5990 9525 -5980
rect 9350 -6010 9495 -5990
rect 9515 -6010 9525 -5990
rect 9350 -6020 9525 -6010
rect 6450 -6415 6465 -6260
rect 6520 -6415 6530 -6260
rect 9435 -6140 9515 -6110
rect 9435 -6295 9445 -6140
rect 9500 -6295 9515 -6140
rect 9280 -6325 9515 -6295
rect 9555 -6140 9635 -5885
rect 9555 -6295 9570 -6140
rect 9625 -6295 9635 -6140
rect 9555 -6310 9635 -6295
rect 9280 -6330 9375 -6325
rect 9280 -6335 9320 -6330
rect 9280 -6360 9290 -6335
rect 9310 -6360 9320 -6335
rect 9280 -6365 9320 -6360
rect 9435 -6350 9515 -6325
rect 9435 -6370 9450 -6350
rect 9490 -6370 9515 -6350
rect 9435 -6380 9515 -6370
rect 6450 -6430 6530 -6415
rect 6175 -6450 6270 -6445
rect 6175 -6455 6215 -6450
rect 6175 -6480 6185 -6455
rect 6205 -6480 6215 -6455
rect 6175 -6485 6215 -6480
rect 6330 -6470 6410 -6445
rect 6330 -6490 6345 -6470
rect 6385 -6490 6410 -6470
rect 6330 -6500 6410 -6490
rect 3005 -6535 3085 -6520
rect 2730 -6555 2825 -6550
rect 2730 -6560 2770 -6555
rect 2730 -6585 2740 -6560
rect 2760 -6585 2770 -6560
rect 2730 -6590 2770 -6585
rect 2885 -6575 2965 -6550
rect 2885 -6595 2900 -6575
rect 2940 -6595 2965 -6575
rect 2885 -6605 2965 -6595
<< viali >>
rect 1565 -1815 1585 -1790
rect 2695 -1785 2715 -1760
rect 4870 -1780 4890 -1755
rect 6000 -1750 6020 -1725
rect 8175 -1745 8195 -1720
rect 9305 -1715 9325 -1690
rect 11480 -1710 11500 -1685
rect 12610 -1680 12630 -1655
rect 12845 -1745 12865 -1725
rect 9540 -1780 9560 -1760
rect 6235 -1815 6255 -1795
rect 2930 -1850 2950 -1830
rect -85 -1885 -65 -1860
rect 195 -1885 240 -1860
rect 505 -1895 525 -1875
rect 665 -1900 750 -1865
rect 1000 -1895 1020 -1870
rect 1280 -1895 1325 -1870
rect 1800 -1880 1820 -1860
rect 130 -2245 160 -2220
rect 220 -2405 240 -2380
rect 365 -2380 385 -2360
rect 630 -2410 650 -2390
rect 2090 -1895 2110 -1875
rect 2250 -1900 2335 -1865
rect 3220 -1850 3240 -1825
rect 3500 -1850 3545 -1825
rect 3810 -1860 3830 -1840
rect 1215 -2255 1245 -2230
rect 1305 -2415 1325 -2390
rect 1855 -2390 1875 -2370
rect 720 -2490 740 -2470
rect 835 -2475 855 -2455
rect -45 -2755 -25 -2730
rect 185 -2755 235 -2730
rect 490 -2740 535 -2710
rect 680 -2750 740 -2710
rect 2215 -2410 2235 -2390
rect 3970 -1865 4055 -1830
rect 4305 -1860 4325 -1835
rect 4585 -1860 4630 -1835
rect 5105 -1845 5125 -1825
rect 3435 -2210 3465 -2185
rect 2985 -2360 3005 -2340
rect 2305 -2490 2325 -2470
rect 3525 -2370 3545 -2345
rect 3670 -2345 3690 -2325
rect 3935 -2375 3955 -2355
rect 5395 -1860 5415 -1840
rect 5555 -1865 5640 -1830
rect 6525 -1815 6545 -1790
rect 6805 -1815 6850 -1790
rect 7115 -1825 7135 -1805
rect 4520 -2220 4550 -2195
rect 4610 -2380 4630 -2355
rect 5160 -2355 5180 -2335
rect 4025 -2455 4045 -2435
rect 4140 -2440 4160 -2420
rect 1040 -2765 1060 -2740
rect 1270 -2765 1320 -2740
rect 1580 -2765 1600 -2740
rect 1795 -2745 1820 -2725
rect 2075 -2740 2120 -2710
rect 2265 -2750 2325 -2710
rect 2710 -2735 2730 -2710
rect 2925 -2715 2950 -2695
rect 3260 -2720 3280 -2695
rect 3490 -2720 3540 -2695
rect 3795 -2705 3840 -2675
rect 3985 -2715 4045 -2675
rect 5520 -2375 5540 -2355
rect 7275 -1830 7360 -1795
rect 7610 -1825 7630 -1800
rect 7890 -1825 7935 -1800
rect 8410 -1810 8430 -1790
rect 6740 -2175 6770 -2150
rect 6290 -2325 6310 -2305
rect 5610 -2455 5630 -2435
rect 6830 -2335 6850 -2310
rect 6975 -2310 6995 -2290
rect 7240 -2340 7260 -2320
rect 8700 -1825 8720 -1805
rect 8860 -1830 8945 -1795
rect 9830 -1780 9850 -1755
rect 10110 -1780 10155 -1755
rect 10420 -1790 10440 -1770
rect 7825 -2185 7855 -2160
rect 7915 -2345 7935 -2320
rect 8465 -2320 8485 -2300
rect 7330 -2420 7350 -2400
rect 7445 -2405 7465 -2385
rect 4345 -2730 4365 -2705
rect 4575 -2730 4625 -2705
rect 4885 -2730 4905 -2705
rect 5100 -2710 5125 -2690
rect 5380 -2705 5425 -2675
rect 5570 -2715 5630 -2675
rect 6015 -2700 6035 -2675
rect 6230 -2680 6255 -2660
rect 6565 -2685 6585 -2660
rect 6795 -2685 6845 -2660
rect 7100 -2670 7145 -2640
rect 7290 -2680 7350 -2640
rect 8825 -2340 8845 -2320
rect 10580 -1795 10665 -1760
rect 10915 -1790 10935 -1765
rect 11195 -1790 11240 -1765
rect 11715 -1775 11735 -1755
rect 10045 -2140 10075 -2115
rect 9595 -2290 9615 -2270
rect 8915 -2420 8935 -2400
rect 10135 -2300 10155 -2275
rect 10280 -2275 10300 -2255
rect 10545 -2305 10565 -2285
rect 12005 -1790 12025 -1770
rect 12165 -1795 12250 -1760
rect 11130 -2150 11160 -2125
rect 11220 -2310 11240 -2285
rect 11770 -2285 11790 -2265
rect 10635 -2385 10655 -2365
rect 10750 -2370 10770 -2350
rect 7650 -2695 7670 -2670
rect 7880 -2695 7930 -2670
rect 8190 -2695 8210 -2670
rect 8405 -2675 8430 -2655
rect 8685 -2670 8730 -2640
rect 8875 -2680 8935 -2640
rect 9320 -2665 9340 -2640
rect 9535 -2645 9560 -2625
rect 9870 -2650 9890 -2625
rect 10100 -2650 10150 -2625
rect 10405 -2635 10450 -2605
rect 10595 -2645 10655 -2605
rect 12130 -2305 12150 -2285
rect 12900 -2255 12920 -2235
rect 12220 -2385 12240 -2365
rect 10955 -2660 10975 -2635
rect 11185 -2660 11235 -2635
rect 11495 -2660 11515 -2635
rect 11710 -2640 11735 -2620
rect 11990 -2635 12035 -2605
rect 12180 -2645 12240 -2605
rect 12625 -2630 12645 -2605
rect 12840 -2610 12865 -2590
rect 130 -2965 150 -2940
rect 948 -2940 968 -2915
rect 3435 -2930 3455 -2905
rect 4253 -2905 4273 -2880
rect 6740 -2895 6760 -2870
rect 7558 -2870 7578 -2845
rect 10045 -2860 10065 -2835
rect 10863 -2835 10883 -2810
rect 365 -3030 385 -3010
rect 945 -3150 965 -3130
rect 3670 -2995 3690 -2975
rect 943 -3535 963 -3510
rect 1655 -3465 1675 -3440
rect 940 -3765 960 -3745
rect 145 -3915 165 -3890
rect 360 -3895 385 -3875
rect 1890 -3530 1910 -3510
rect 2473 -3440 2493 -3415
rect 4250 -3115 4270 -3095
rect 6975 -2960 6995 -2940
rect 4248 -3500 4268 -3475
rect 4960 -3430 4980 -3405
rect 2735 -3735 2755 -3710
rect 2880 -3800 2930 -3775
rect 2468 -4035 2488 -4010
rect 80 -4225 100 -4200
rect 898 -4200 918 -4175
rect 315 -4290 335 -4270
rect 895 -4410 915 -4390
rect 1670 -4415 1690 -4390
rect 1885 -4395 1910 -4375
rect 4245 -3730 4265 -3710
rect 3450 -3880 3470 -3855
rect 3665 -3860 3690 -3840
rect 5195 -3495 5215 -3475
rect 5778 -3405 5798 -3380
rect 7555 -3080 7575 -3060
rect 10280 -2925 10300 -2905
rect 7553 -3465 7573 -3440
rect 8265 -3395 8285 -3370
rect 6065 -3700 6085 -3675
rect 6210 -3765 6260 -3740
rect 5773 -4000 5793 -3975
rect 3385 -4190 3405 -4165
rect 4203 -4165 4223 -4140
rect 3620 -4255 3640 -4235
rect 893 -4795 913 -4770
rect 2665 -4765 2685 -4740
rect 2825 -4775 2865 -4755
rect 890 -5025 910 -5005
rect 95 -5175 115 -5150
rect 310 -5155 335 -5135
rect 4200 -4375 4220 -4355
rect 4975 -4380 4995 -4355
rect 5190 -4360 5215 -4340
rect 7550 -3695 7570 -3675
rect 6755 -3845 6775 -3820
rect 6970 -3825 6995 -3805
rect 8500 -3460 8520 -3440
rect 9083 -3370 9103 -3345
rect 10860 -3045 10880 -3025
rect 13650 -3090 13670 -3065
rect 13220 -3130 13240 -3105
rect 13795 -3155 13845 -3130
rect 13365 -3195 13415 -3170
rect 10858 -3430 10878 -3405
rect 11570 -3360 11590 -3335
rect 9380 -3665 9400 -3640
rect 9525 -3730 9575 -3705
rect 9078 -3965 9098 -3940
rect 6690 -4155 6710 -4130
rect 7508 -4130 7528 -4105
rect 6925 -4220 6945 -4200
rect 4198 -4760 4218 -4735
rect 5995 -4730 6015 -4705
rect 6155 -4740 6195 -4720
rect 4195 -4990 4215 -4970
rect 3400 -5140 3420 -5115
rect 3615 -5120 3640 -5100
rect 7505 -4340 7525 -4320
rect 8280 -4345 8300 -4320
rect 8495 -4325 8520 -4305
rect 10855 -3660 10875 -3640
rect 10060 -3810 10080 -3785
rect 10275 -3790 10300 -3770
rect 11805 -3425 11825 -3405
rect 12388 -3335 12408 -3310
rect 12383 -3930 12403 -3905
rect 9995 -4120 10015 -4095
rect 10813 -4095 10833 -4070
rect 10230 -4185 10250 -4165
rect 7503 -4725 7523 -4700
rect 9310 -4695 9330 -4670
rect 9470 -4705 9510 -4685
rect 2810 -5555 2830 -5530
rect 2955 -5620 3005 -5595
rect 7500 -4955 7520 -4935
rect 6705 -5105 6725 -5080
rect 6920 -5085 6945 -5065
rect 10810 -4305 10830 -4285
rect 11585 -4310 11605 -4285
rect 11800 -4290 11825 -4270
rect 13580 -4120 13600 -4095
rect 13150 -4160 13170 -4135
rect 13740 -4130 13780 -4110
rect 13310 -4170 13350 -4150
rect 10808 -4690 10828 -4665
rect 6255 -5450 6275 -5425
rect 10805 -4920 10825 -4900
rect 10010 -5070 10030 -5045
rect 10225 -5050 10250 -5030
rect 9360 -5330 9380 -5305
rect 9505 -5395 9555 -5370
rect 6400 -5515 6450 -5490
rect 9290 -6360 9310 -6335
rect 9450 -6370 9490 -6350
rect 6185 -6480 6205 -6455
rect 6345 -6490 6385 -6470
rect 2740 -6585 2760 -6560
rect 2900 -6595 2940 -6575
<< metal1 >>
rect 12605 -1655 12635 -1645
rect 9300 -1690 9330 -1680
rect 5995 -1725 6025 -1715
rect 2690 -1760 2720 -1750
rect 1560 -1790 1590 -1780
rect 1560 -1815 1565 -1790
rect 1585 -1815 1590 -1790
rect -160 -1855 400 -1845
rect 1560 -1855 1590 -1815
rect 2690 -1785 2695 -1760
rect 2715 -1785 2720 -1760
rect 2690 -1825 2720 -1785
rect 4865 -1755 4895 -1745
rect 4865 -1780 4870 -1755
rect 4890 -1780 4895 -1755
rect 3090 -1815 3705 -1810
rect 2770 -1820 3705 -1815
rect 4865 -1820 4895 -1780
rect 5995 -1750 6000 -1725
rect 6020 -1750 6025 -1725
rect 5995 -1790 6025 -1750
rect 8170 -1720 8200 -1710
rect 8170 -1745 8175 -1720
rect 8195 -1745 8200 -1720
rect 6450 -1780 7010 -1775
rect 6075 -1785 7010 -1780
rect 8170 -1785 8200 -1745
rect 9300 -1715 9305 -1690
rect 9325 -1715 9330 -1690
rect 9300 -1755 9330 -1715
rect 11475 -1685 11505 -1675
rect 11475 -1710 11480 -1685
rect 11500 -1710 11505 -1685
rect 9755 -1745 10315 -1740
rect 9380 -1750 10315 -1745
rect 11475 -1750 11505 -1710
rect 12605 -1680 12610 -1655
rect 12630 -1680 12635 -1655
rect 12605 -1720 12635 -1680
rect 12685 -1720 13245 -1710
rect 12500 -1725 13245 -1720
rect 11555 -1745 11825 -1740
rect 12500 -1745 12845 -1725
rect 12865 -1745 13245 -1725
rect 11555 -1750 11885 -1745
rect 12500 -1750 13245 -1745
rect 9380 -1755 13245 -1750
rect 9195 -1760 9830 -1755
rect 8250 -1780 8520 -1775
rect 9195 -1780 9540 -1760
rect 9560 -1780 9830 -1760
rect 9850 -1780 10110 -1755
rect 10155 -1760 11715 -1755
rect 10155 -1770 10580 -1760
rect 10155 -1780 10420 -1770
rect 8250 -1785 8580 -1780
rect 9195 -1785 10420 -1780
rect 6075 -1790 10315 -1785
rect 10370 -1790 10420 -1785
rect 10440 -1790 10580 -1770
rect 5890 -1795 6525 -1790
rect 4945 -1815 5215 -1810
rect 5890 -1815 6235 -1795
rect 6255 -1815 6525 -1795
rect 6545 -1815 6805 -1790
rect 6850 -1795 8410 -1790
rect 6850 -1805 7275 -1795
rect 6850 -1815 7115 -1805
rect 4945 -1820 5275 -1815
rect 5890 -1820 7115 -1815
rect 2770 -1825 7010 -1820
rect 7065 -1825 7115 -1820
rect 7135 -1825 7275 -1805
rect 2585 -1830 3220 -1825
rect 1640 -1850 1910 -1845
rect 2585 -1850 2930 -1830
rect 2950 -1850 3220 -1830
rect 3240 -1850 3500 -1825
rect 3545 -1830 5105 -1825
rect 3545 -1840 3970 -1830
rect 3545 -1850 3810 -1840
rect 1640 -1855 1970 -1850
rect 2585 -1855 3810 -1850
rect -160 -1860 3705 -1855
rect 3760 -1860 3810 -1855
rect 3830 -1860 3970 -1840
rect -160 -1885 -85 -1860
rect -65 -1885 195 -1860
rect 240 -1865 1800 -1860
rect 240 -1875 665 -1865
rect 240 -1885 505 -1875
rect -160 -1890 505 -1885
rect -160 -1895 400 -1890
rect 455 -1895 505 -1890
rect 525 -1895 665 -1875
rect -160 -2930 -135 -1895
rect 455 -1900 665 -1895
rect 750 -1870 1800 -1865
rect 750 -1895 1000 -1870
rect 1020 -1895 1280 -1870
rect 1325 -1880 1800 -1870
rect 1820 -1865 2770 -1860
rect 1820 -1875 2250 -1865
rect 1820 -1880 2090 -1875
rect 1325 -1890 2090 -1880
rect 1325 -1895 1640 -1890
rect 750 -1900 1640 -1895
rect 455 -1905 1640 -1900
rect 2045 -1895 2090 -1890
rect 2110 -1895 2250 -1875
rect 2045 -1900 2250 -1895
rect 2335 -1875 2770 -1865
rect 3760 -1865 3970 -1860
rect 4055 -1835 5105 -1830
rect 4055 -1860 4305 -1835
rect 4325 -1860 4585 -1835
rect 4630 -1845 5105 -1835
rect 5125 -1830 6075 -1825
rect 5125 -1840 5555 -1830
rect 5125 -1845 5395 -1840
rect 4630 -1855 5395 -1845
rect 4630 -1860 4945 -1855
rect 4055 -1865 4945 -1860
rect 3760 -1870 4945 -1865
rect 5350 -1860 5395 -1855
rect 5415 -1860 5555 -1840
rect 5350 -1865 5555 -1860
rect 5640 -1840 6075 -1830
rect 7065 -1830 7275 -1825
rect 7360 -1800 8410 -1795
rect 7360 -1825 7610 -1800
rect 7630 -1825 7890 -1800
rect 7935 -1810 8410 -1800
rect 8430 -1795 9380 -1790
rect 8430 -1805 8860 -1795
rect 8430 -1810 8700 -1805
rect 7935 -1820 8700 -1810
rect 7935 -1825 8250 -1820
rect 7360 -1830 8250 -1825
rect 7065 -1835 8250 -1830
rect 8655 -1825 8700 -1820
rect 8720 -1825 8860 -1805
rect 8655 -1830 8860 -1825
rect 8945 -1805 9380 -1795
rect 10370 -1795 10580 -1790
rect 10665 -1765 11715 -1760
rect 10665 -1790 10915 -1765
rect 10935 -1790 11195 -1765
rect 11240 -1775 11715 -1765
rect 11735 -1760 12685 -1755
rect 11735 -1770 12165 -1760
rect 11735 -1775 12005 -1770
rect 11240 -1785 12005 -1775
rect 11240 -1790 11555 -1785
rect 10665 -1795 11555 -1790
rect 10370 -1800 11555 -1795
rect 11960 -1790 12005 -1785
rect 12025 -1790 12165 -1770
rect 11960 -1795 12165 -1790
rect 12250 -1770 12685 -1760
rect 12250 -1780 12525 -1770
rect 12250 -1795 12515 -1780
rect 8945 -1815 9220 -1805
rect 10370 -1810 10895 -1800
rect 11960 -1810 12515 -1795
rect 8945 -1830 9210 -1815
rect 5640 -1850 5915 -1840
rect 7065 -1845 7590 -1835
rect 8655 -1845 9210 -1830
rect 5640 -1865 5905 -1850
rect 2335 -1885 2610 -1875
rect 3760 -1880 4285 -1870
rect 5350 -1880 5905 -1865
rect 2335 -1900 2600 -1885
rect 455 -1915 980 -1905
rect 2045 -1915 2600 -1900
rect 10035 -2115 10085 -2105
rect 10035 -2140 10045 -2115
rect 10075 -2140 10085 -2115
rect 6730 -2150 6780 -2140
rect 10035 -2150 10085 -2140
rect 11120 -2125 11170 -2115
rect 11120 -2150 11130 -2125
rect 11160 -2150 11170 -2125
rect 6730 -2175 6740 -2150
rect 6770 -2175 6780 -2150
rect 3425 -2185 3475 -2175
rect 6730 -2185 6780 -2175
rect 7815 -2160 7865 -2150
rect 11120 -2160 11170 -2150
rect 7815 -2185 7825 -2160
rect 7855 -2185 7865 -2160
rect 3425 -2210 3435 -2185
rect 3465 -2210 3475 -2185
rect 120 -2220 170 -2210
rect 3425 -2220 3475 -2210
rect 4510 -2195 4560 -2185
rect 7815 -2195 7865 -2185
rect 4510 -2220 4520 -2195
rect 4550 -2220 4560 -2195
rect 120 -2245 130 -2220
rect 160 -2245 170 -2220
rect 120 -2255 170 -2245
rect 1205 -2230 1255 -2220
rect 4510 -2230 4560 -2220
rect 12890 -2230 12930 -2225
rect 1205 -2255 1215 -2230
rect 1245 -2255 1255 -2230
rect 1205 -2265 1255 -2255
rect 10270 -2250 10310 -2245
rect 9585 -2265 9625 -2260
rect 6965 -2285 7005 -2280
rect 6280 -2300 6320 -2295
rect 3660 -2320 3700 -2315
rect 2975 -2335 3015 -2330
rect 355 -2355 395 -2350
rect 210 -2380 250 -2370
rect 210 -2405 220 -2380
rect 240 -2405 250 -2380
rect 355 -2385 360 -2355
rect 390 -2385 395 -2355
rect 1845 -2365 1885 -2360
rect 355 -2390 395 -2385
rect 620 -2390 660 -2385
rect 210 -2415 250 -2405
rect 620 -2410 630 -2390
rect 650 -2410 660 -2390
rect 620 -2415 660 -2410
rect 1295 -2390 1335 -2380
rect 1295 -2415 1305 -2390
rect 1325 -2415 1335 -2390
rect 1845 -2395 1850 -2365
rect 1880 -2395 1885 -2365
rect 2975 -2365 2980 -2335
rect 3010 -2365 3015 -2335
rect 2975 -2370 3015 -2365
rect 3515 -2345 3555 -2335
rect 3515 -2370 3525 -2345
rect 3545 -2370 3555 -2345
rect 3660 -2350 3665 -2320
rect 3695 -2350 3700 -2320
rect 5150 -2330 5190 -2325
rect 3660 -2355 3700 -2350
rect 3925 -2355 3965 -2350
rect 3515 -2380 3555 -2370
rect 3925 -2375 3935 -2355
rect 3955 -2375 3965 -2355
rect 3925 -2380 3965 -2375
rect 4600 -2355 4640 -2345
rect 4600 -2380 4610 -2355
rect 4630 -2380 4640 -2355
rect 5150 -2360 5155 -2330
rect 5185 -2360 5190 -2330
rect 6280 -2330 6285 -2300
rect 6315 -2330 6320 -2300
rect 6280 -2335 6320 -2330
rect 6820 -2310 6860 -2300
rect 6820 -2335 6830 -2310
rect 6850 -2335 6860 -2310
rect 6965 -2315 6970 -2285
rect 7000 -2315 7005 -2285
rect 8455 -2295 8495 -2290
rect 6965 -2320 7005 -2315
rect 7230 -2320 7270 -2315
rect 6820 -2345 6860 -2335
rect 7230 -2340 7240 -2320
rect 7260 -2340 7270 -2320
rect 7230 -2345 7270 -2340
rect 7905 -2320 7945 -2310
rect 7905 -2345 7915 -2320
rect 7935 -2345 7945 -2320
rect 8455 -2325 8460 -2295
rect 8490 -2325 8495 -2295
rect 9585 -2295 9590 -2265
rect 9620 -2295 9625 -2265
rect 9585 -2300 9625 -2295
rect 10125 -2275 10165 -2265
rect 10125 -2300 10135 -2275
rect 10155 -2300 10165 -2275
rect 10270 -2280 10275 -2250
rect 10305 -2280 10310 -2250
rect 11760 -2260 11800 -2255
rect 10270 -2285 10310 -2280
rect 10535 -2285 10575 -2280
rect 10125 -2310 10165 -2300
rect 10535 -2305 10545 -2285
rect 10565 -2305 10575 -2285
rect 10535 -2310 10575 -2305
rect 11210 -2285 11250 -2275
rect 11210 -2310 11220 -2285
rect 11240 -2310 11250 -2285
rect 11760 -2290 11765 -2260
rect 11795 -2290 11800 -2260
rect 12890 -2260 12895 -2230
rect 12925 -2260 12930 -2230
rect 12890 -2265 12930 -2260
rect 11760 -2295 11800 -2290
rect 12120 -2285 12160 -2280
rect 12120 -2305 12130 -2285
rect 12150 -2305 12160 -2285
rect 12120 -2310 12160 -2305
rect 8455 -2330 8495 -2325
rect 8815 -2320 8855 -2315
rect 11210 -2320 11250 -2310
rect 8815 -2340 8825 -2320
rect 8845 -2340 8855 -2320
rect 8815 -2345 8855 -2340
rect 10740 -2345 10780 -2340
rect 5150 -2365 5190 -2360
rect 5510 -2355 5550 -2350
rect 7905 -2355 7945 -2345
rect 5510 -2375 5520 -2355
rect 5540 -2375 5550 -2355
rect 10625 -2365 10665 -2360
rect 5510 -2380 5550 -2375
rect 7435 -2380 7475 -2375
rect 1845 -2400 1885 -2395
rect 2205 -2390 2245 -2385
rect 4600 -2390 4640 -2380
rect 2205 -2410 2215 -2390
rect 2235 -2410 2245 -2390
rect 7320 -2400 7360 -2395
rect 2205 -2415 2245 -2410
rect 4130 -2415 4170 -2410
rect 1295 -2425 1335 -2415
rect 4015 -2435 4055 -2430
rect 825 -2450 865 -2445
rect 710 -2470 750 -2465
rect 710 -2490 720 -2470
rect 740 -2490 750 -2470
rect 825 -2480 830 -2450
rect 860 -2480 865 -2450
rect 4015 -2455 4025 -2435
rect 4045 -2455 4055 -2435
rect 4130 -2445 4135 -2415
rect 4165 -2445 4170 -2415
rect 7320 -2420 7330 -2400
rect 7350 -2420 7360 -2400
rect 7435 -2410 7440 -2380
rect 7470 -2410 7475 -2380
rect 10625 -2385 10635 -2365
rect 10655 -2385 10665 -2365
rect 10740 -2375 10745 -2345
rect 10775 -2375 10780 -2345
rect 10740 -2380 10780 -2375
rect 12210 -2365 12250 -2360
rect 10625 -2390 10665 -2385
rect 12210 -2385 12220 -2365
rect 12240 -2385 12250 -2365
rect 12210 -2390 12250 -2385
rect 7435 -2415 7475 -2410
rect 8905 -2400 8945 -2395
rect 7320 -2425 7360 -2420
rect 8905 -2420 8915 -2400
rect 8935 -2420 8945 -2400
rect 8905 -2425 8945 -2420
rect 4130 -2450 4170 -2445
rect 5600 -2435 5640 -2430
rect 4015 -2460 4055 -2455
rect 5600 -2455 5610 -2435
rect 5630 -2455 5640 -2435
rect 5600 -2460 5640 -2455
rect 825 -2485 865 -2480
rect 2295 -2470 2335 -2465
rect 710 -2495 750 -2490
rect 2295 -2490 2305 -2470
rect 2325 -2490 2335 -2470
rect 2295 -2495 2335 -2490
rect 12725 -2590 12955 -2580
rect 10395 -2605 10460 -2595
rect 10370 -2615 10405 -2605
rect 9420 -2625 10405 -2615
rect 7090 -2640 7155 -2630
rect 7065 -2650 7100 -2640
rect 6115 -2660 7100 -2650
rect 3785 -2675 3850 -2665
rect 3760 -2685 3795 -2675
rect 2810 -2695 3795 -2685
rect 480 -2710 545 -2700
rect 455 -2720 490 -2710
rect -55 -2730 490 -2720
rect -55 -2755 -45 -2730
rect -25 -2755 185 -2730
rect 235 -2740 490 -2730
rect 535 -2740 545 -2710
rect 235 -2750 545 -2740
rect 600 -2710 875 -2695
rect 600 -2750 680 -2710
rect 740 -2735 875 -2710
rect 2045 -2700 2075 -2695
rect 2185 -2700 2700 -2695
rect 2810 -2700 2925 -2695
rect 2045 -2710 2130 -2700
rect 2045 -2715 2075 -2710
rect 955 -2730 1010 -2720
rect 1680 -2725 2075 -2715
rect 1680 -2730 1795 -2725
rect 955 -2735 1795 -2730
rect 740 -2740 1795 -2735
rect 740 -2750 1040 -2740
rect 235 -2755 485 -2750
rect 600 -2755 1040 -2750
rect -55 -2765 400 -2755
rect 870 -2765 1040 -2755
rect 1060 -2765 1270 -2740
rect 1320 -2765 1580 -2740
rect 1600 -2745 1795 -2740
rect 1820 -2740 2075 -2725
rect 2120 -2740 2130 -2710
rect 1820 -2745 2130 -2740
rect 1600 -2750 2130 -2745
rect 2185 -2710 2925 -2700
rect 2185 -2750 2265 -2710
rect 2325 -2735 2710 -2710
rect 2730 -2715 2925 -2710
rect 2950 -2715 3260 -2695
rect 2730 -2720 3260 -2715
rect 3280 -2720 3490 -2695
rect 3540 -2705 3795 -2695
rect 3840 -2705 3850 -2675
rect 3540 -2715 3850 -2705
rect 3905 -2675 4180 -2660
rect 3905 -2715 3985 -2675
rect 4045 -2700 4180 -2675
rect 5350 -2665 5380 -2660
rect 5490 -2665 6005 -2660
rect 6115 -2665 6230 -2660
rect 5350 -2675 5435 -2665
rect 5350 -2680 5380 -2675
rect 4260 -2695 4315 -2685
rect 4985 -2690 5380 -2680
rect 4985 -2695 5100 -2690
rect 4260 -2700 5100 -2695
rect 4045 -2705 5100 -2700
rect 4045 -2715 4345 -2705
rect 3540 -2720 3790 -2715
rect 3905 -2720 4345 -2715
rect 2730 -2735 2810 -2720
rect 3250 -2730 3705 -2720
rect 4175 -2730 4345 -2720
rect 4365 -2730 4575 -2705
rect 4625 -2730 4885 -2705
rect 4905 -2710 5100 -2705
rect 5125 -2705 5380 -2690
rect 5425 -2705 5435 -2675
rect 5125 -2710 5435 -2705
rect 4905 -2715 5435 -2710
rect 5490 -2675 6230 -2665
rect 5490 -2715 5570 -2675
rect 5630 -2700 6015 -2675
rect 6035 -2680 6230 -2675
rect 6255 -2680 6565 -2660
rect 6035 -2685 6565 -2680
rect 6585 -2685 6795 -2660
rect 6845 -2670 7100 -2660
rect 7145 -2670 7155 -2640
rect 6845 -2680 7155 -2670
rect 7210 -2640 7485 -2625
rect 7210 -2680 7290 -2640
rect 7350 -2665 7485 -2640
rect 8655 -2630 8685 -2625
rect 8795 -2630 9310 -2625
rect 9420 -2630 9535 -2625
rect 8655 -2640 8740 -2630
rect 8655 -2645 8685 -2640
rect 7565 -2660 7620 -2650
rect 8290 -2655 8685 -2645
rect 8290 -2660 8405 -2655
rect 7565 -2665 8405 -2660
rect 7350 -2670 8405 -2665
rect 7350 -2680 7650 -2670
rect 6845 -2685 7095 -2680
rect 7210 -2685 7650 -2680
rect 6035 -2700 6115 -2685
rect 6555 -2695 7010 -2685
rect 7480 -2695 7650 -2685
rect 7670 -2695 7880 -2670
rect 7930 -2695 8190 -2670
rect 8210 -2675 8405 -2670
rect 8430 -2670 8685 -2655
rect 8730 -2670 8740 -2640
rect 8430 -2675 8740 -2670
rect 8210 -2680 8740 -2675
rect 8795 -2640 9535 -2630
rect 8795 -2680 8875 -2640
rect 8935 -2665 9320 -2640
rect 9340 -2645 9535 -2640
rect 9560 -2645 9870 -2625
rect 9340 -2650 9870 -2645
rect 9890 -2650 10100 -2625
rect 10150 -2635 10405 -2625
rect 10450 -2635 10460 -2605
rect 10150 -2645 10460 -2635
rect 10515 -2605 10790 -2590
rect 10515 -2645 10595 -2605
rect 10655 -2630 10790 -2605
rect 11960 -2595 11990 -2590
rect 12100 -2595 12615 -2590
rect 12725 -2595 12840 -2590
rect 11960 -2605 12045 -2595
rect 11960 -2610 11990 -2605
rect 10870 -2625 10925 -2615
rect 11595 -2620 11990 -2610
rect 11595 -2625 11710 -2620
rect 10870 -2630 11710 -2625
rect 10655 -2635 11710 -2630
rect 10655 -2645 10955 -2635
rect 10150 -2650 10400 -2645
rect 10515 -2650 10955 -2645
rect 9340 -2665 9420 -2650
rect 9860 -2660 10315 -2650
rect 10785 -2660 10955 -2650
rect 10975 -2660 11185 -2635
rect 11235 -2660 11495 -2635
rect 11515 -2640 11710 -2635
rect 11735 -2635 11990 -2620
rect 12035 -2635 12045 -2605
rect 11735 -2640 12045 -2635
rect 11515 -2645 12045 -2640
rect 12100 -2605 12840 -2595
rect 12100 -2645 12180 -2605
rect 12240 -2630 12625 -2605
rect 12645 -2610 12840 -2605
rect 12865 -2610 12955 -2590
rect 12645 -2615 12955 -2610
rect 12645 -2630 12725 -2615
rect 12240 -2640 12725 -2630
rect 12240 -2645 12615 -2640
rect 11515 -2660 11595 -2645
rect 11960 -2660 11990 -2645
rect 12100 -2650 12615 -2645
rect 8935 -2675 9420 -2665
rect 10785 -2665 11595 -2660
rect 10785 -2670 10925 -2665
rect 10945 -2670 11595 -2665
rect 10870 -2675 10925 -2670
rect 8935 -2680 9310 -2675
rect 8210 -2695 8290 -2680
rect 8655 -2695 8685 -2680
rect 8795 -2685 9310 -2680
rect 5630 -2710 6115 -2700
rect 7480 -2700 8290 -2695
rect 7480 -2705 7620 -2700
rect 7640 -2705 8290 -2700
rect 7565 -2710 7620 -2705
rect 5630 -2715 6005 -2710
rect 4905 -2730 4985 -2715
rect 5350 -2730 5380 -2715
rect 5490 -2720 6005 -2715
rect 2325 -2745 2810 -2735
rect 4175 -2735 4985 -2730
rect 4175 -2740 4315 -2735
rect 4335 -2740 4985 -2735
rect 4260 -2745 4315 -2740
rect 2325 -2750 2700 -2745
rect 1600 -2765 1680 -2750
rect 2045 -2765 2075 -2750
rect 2185 -2755 2700 -2750
rect 870 -2770 1680 -2765
rect 870 -2775 1010 -2770
rect 1030 -2775 1680 -2770
rect 10545 -2775 11595 -2745
rect 955 -2780 1010 -2775
rect 7240 -2810 8290 -2780
rect 3935 -2845 4985 -2815
rect 630 -2880 1680 -2850
rect -160 -2935 155 -2930
rect -370 -2940 155 -2935
rect -370 -2965 130 -2940
rect 150 -2965 155 -2940
rect -370 -2970 155 -2965
rect -370 -5625 -295 -2970
rect -160 -2975 155 -2970
rect 125 -3005 155 -2975
rect 205 -3000 475 -2995
rect 630 -3000 655 -2880
rect 205 -3005 655 -3000
rect 125 -3010 655 -3005
rect 125 -3030 365 -3010
rect 385 -3030 655 -3010
rect 125 -3040 655 -3030
rect 125 -3055 205 -3040
rect 125 -3095 185 -3055
rect 840 -3460 870 -2880
rect 945 -2905 970 -2880
rect 943 -2915 973 -2905
rect 943 -2940 948 -2915
rect 968 -2940 973 -2915
rect 943 -2970 973 -2940
rect 935 -3125 975 -3120
rect 935 -3155 940 -3125
rect 970 -3155 975 -3125
rect 935 -3160 975 -3155
rect 1650 -3250 1680 -2880
rect 3430 -2905 3460 -2895
rect 3430 -2930 3435 -2905
rect 3455 -2930 3460 -2905
rect 3430 -2970 3460 -2930
rect 3510 -2965 3780 -2960
rect 3935 -2965 3960 -2845
rect 3510 -2970 3960 -2965
rect 3430 -2975 3960 -2970
rect 3430 -2995 3670 -2975
rect 3690 -2995 3960 -2975
rect 3430 -3005 3960 -2995
rect 3430 -3020 3510 -3005
rect 3430 -3250 3460 -3020
rect 1650 -3280 3460 -3250
rect 1650 -3440 1680 -3280
rect 2470 -3405 2495 -3280
rect 840 -3475 965 -3460
rect 245 -3875 517 -3865
rect -140 -3890 360 -3875
rect -140 -3915 145 -3890
rect 165 -3895 360 -3890
rect 385 -3895 517 -3875
rect 165 -3900 517 -3895
rect 165 -3915 275 -3900
rect -140 -3935 275 -3915
rect -140 -5135 -95 -3935
rect 840 -4120 870 -3475
rect 940 -3500 965 -3475
rect 1650 -3465 1655 -3440
rect 1675 -3465 1680 -3440
rect 938 -3510 968 -3500
rect 1650 -3505 1680 -3465
rect 2468 -3415 2498 -3405
rect 2468 -3440 2473 -3415
rect 2493 -3440 2498 -3415
rect 2468 -3470 2498 -3440
rect 1730 -3500 2000 -3495
rect 1730 -3505 2190 -3500
rect 938 -3535 943 -3510
rect 963 -3535 968 -3510
rect 1590 -3510 2190 -3505
rect 1590 -3530 1890 -3510
rect 1910 -3530 2190 -3510
rect 1590 -3535 2190 -3530
rect 938 -3565 968 -3535
rect 1548 -3540 2190 -3535
rect 1548 -3555 1730 -3540
rect 1548 -3595 1710 -3555
rect 930 -3740 970 -3735
rect 930 -3770 935 -3740
rect 965 -3770 970 -3740
rect 930 -3775 970 -3770
rect 2165 -3935 2190 -3540
rect 2730 -3710 2760 -3700
rect 2730 -3735 2735 -3710
rect 2755 -3735 2760 -3710
rect 2730 -3775 2760 -3735
rect 3030 -3765 3070 -3280
rect 2810 -3775 3070 -3765
rect 2670 -3800 2880 -3775
rect 2930 -3800 3070 -3775
rect 2670 -3805 3070 -3800
rect 2628 -3810 3070 -3805
rect 4145 -3425 4175 -2845
rect 4250 -2870 4275 -2845
rect 4248 -2880 4278 -2870
rect 4248 -2905 4253 -2880
rect 4273 -2905 4278 -2880
rect 4248 -2935 4278 -2905
rect 4240 -3090 4280 -3085
rect 4240 -3120 4245 -3090
rect 4275 -3120 4280 -3090
rect 4240 -3125 4280 -3120
rect 4955 -3215 4985 -2845
rect 6735 -2870 6765 -2860
rect 6735 -2895 6740 -2870
rect 6760 -2895 6765 -2870
rect 6735 -2935 6765 -2895
rect 6815 -2930 7085 -2925
rect 7240 -2930 7265 -2810
rect 6815 -2935 7265 -2930
rect 6735 -2940 7265 -2935
rect 6735 -2960 6975 -2940
rect 6995 -2960 7265 -2940
rect 6735 -2970 7265 -2960
rect 6735 -2985 6815 -2970
rect 6735 -3215 6765 -2985
rect 4955 -3245 6765 -3215
rect 4955 -3405 4985 -3245
rect 5775 -3370 5800 -3245
rect 4145 -3440 4270 -3425
rect 2628 -3825 2810 -3810
rect 2628 -3865 2790 -3825
rect 3550 -3840 3822 -3830
rect 3165 -3855 3665 -3840
rect 3165 -3880 3450 -3855
rect 3470 -3860 3665 -3855
rect 3690 -3860 3822 -3840
rect 3470 -3865 3822 -3860
rect 3470 -3880 3580 -3865
rect 3165 -3900 3580 -3880
rect 2165 -3960 2490 -3935
rect 2465 -4000 2490 -3960
rect 2463 -4010 2493 -4000
rect 2463 -4035 2468 -4010
rect 2488 -4035 2493 -4010
rect 2463 -4065 2493 -4035
rect 595 -4140 920 -4120
rect 75 -4200 105 -4190
rect 75 -4225 80 -4200
rect 100 -4225 105 -4200
rect 75 -4265 105 -4225
rect 155 -4260 425 -4255
rect 595 -4260 625 -4140
rect 155 -4265 625 -4260
rect 15 -4270 625 -4265
rect 15 -4290 315 -4270
rect 335 -4290 625 -4270
rect 15 -4295 625 -4290
rect -27 -4300 625 -4295
rect -27 -4315 155 -4300
rect -27 -4355 135 -4315
rect 720 -4635 755 -4140
rect 895 -4165 920 -4140
rect 893 -4175 923 -4165
rect 893 -4200 898 -4175
rect 918 -4200 923 -4175
rect 893 -4230 923 -4200
rect 1770 -4375 2042 -4365
rect 885 -4385 925 -4380
rect 885 -4415 890 -4385
rect 920 -4415 925 -4385
rect 885 -4420 925 -4415
rect 1550 -4390 1885 -4375
rect 1550 -4415 1670 -4390
rect 1690 -4395 1885 -4390
rect 1910 -4395 2042 -4375
rect 1690 -4400 2042 -4395
rect 1690 -4415 1800 -4400
rect 1550 -4435 1800 -4415
rect 720 -4660 915 -4635
rect 890 -4760 915 -4660
rect 888 -4770 918 -4760
rect 888 -4795 893 -4770
rect 913 -4795 918 -4770
rect 888 -4825 918 -4795
rect 880 -5000 920 -4995
rect 880 -5030 885 -5000
rect 915 -5030 920 -5000
rect 880 -5035 920 -5030
rect 195 -5135 475 -5125
rect -140 -5150 310 -5135
rect -140 -5175 95 -5150
rect 115 -5155 310 -5150
rect 335 -5155 475 -5135
rect 115 -5160 475 -5155
rect 115 -5175 225 -5160
rect -140 -5195 225 -5175
rect 440 -5215 475 -5160
rect 1550 -5215 1580 -4435
rect 2620 -4740 2750 -4725
rect 2620 -4765 2665 -4740
rect 2685 -4755 3010 -4740
rect 2685 -4765 2825 -4755
rect 2620 -4775 2825 -4765
rect 2865 -4775 3010 -4755
rect 2620 -4785 3010 -4775
rect 2620 -5215 2655 -4785
rect 3165 -5100 3210 -3900
rect 4145 -4085 4175 -3440
rect 4245 -3465 4270 -3440
rect 4955 -3430 4960 -3405
rect 4980 -3430 4985 -3405
rect 4243 -3475 4273 -3465
rect 4955 -3470 4985 -3430
rect 5773 -3380 5803 -3370
rect 5773 -3405 5778 -3380
rect 5798 -3405 5803 -3380
rect 5773 -3435 5803 -3405
rect 5035 -3465 5305 -3460
rect 5035 -3470 5495 -3465
rect 4243 -3500 4248 -3475
rect 4268 -3500 4273 -3475
rect 4895 -3475 5495 -3470
rect 4895 -3495 5195 -3475
rect 5215 -3495 5495 -3475
rect 4895 -3500 5495 -3495
rect 4243 -3530 4273 -3500
rect 4853 -3505 5495 -3500
rect 4853 -3520 5035 -3505
rect 4853 -3560 5015 -3520
rect 4235 -3705 4275 -3700
rect 4235 -3735 4240 -3705
rect 4270 -3735 4275 -3705
rect 4235 -3740 4275 -3735
rect 5470 -3900 5495 -3505
rect 6060 -3675 6090 -3665
rect 6060 -3700 6065 -3675
rect 6085 -3700 6090 -3675
rect 6060 -3740 6090 -3700
rect 6365 -3730 6400 -3245
rect 6140 -3740 6400 -3730
rect 6000 -3765 6210 -3740
rect 6260 -3765 6400 -3740
rect 6000 -3770 6400 -3765
rect 5958 -3775 6400 -3770
rect 7450 -3390 7480 -2810
rect 7555 -2835 7580 -2810
rect 7553 -2845 7583 -2835
rect 7553 -2870 7558 -2845
rect 7578 -2870 7583 -2845
rect 7553 -2900 7583 -2870
rect 7545 -3055 7585 -3050
rect 7545 -3085 7550 -3055
rect 7580 -3085 7585 -3055
rect 7545 -3090 7585 -3085
rect 8260 -3180 8290 -2810
rect 10040 -2835 10070 -2825
rect 10040 -2860 10045 -2835
rect 10065 -2860 10070 -2835
rect 10040 -2900 10070 -2860
rect 10120 -2895 10390 -2890
rect 10545 -2895 10570 -2775
rect 10120 -2900 10570 -2895
rect 10040 -2905 10570 -2900
rect 10040 -2925 10280 -2905
rect 10300 -2925 10570 -2905
rect 10040 -2935 10570 -2925
rect 10040 -2950 10120 -2935
rect 10040 -3180 10070 -2950
rect 8260 -3210 10070 -3180
rect 8260 -3370 8290 -3210
rect 9080 -3335 9105 -3210
rect 7450 -3405 7575 -3390
rect 5958 -3790 6140 -3775
rect 5958 -3830 6120 -3790
rect 6855 -3805 7127 -3795
rect 6470 -3820 6970 -3805
rect 6470 -3845 6755 -3820
rect 6775 -3825 6970 -3820
rect 6995 -3825 7127 -3805
rect 6775 -3830 7127 -3825
rect 6775 -3845 6885 -3830
rect 6470 -3865 6885 -3845
rect 5470 -3925 5795 -3900
rect 5770 -3965 5795 -3925
rect 5768 -3975 5798 -3965
rect 5768 -4000 5773 -3975
rect 5793 -4000 5798 -3975
rect 5768 -4030 5798 -4000
rect 3900 -4105 4225 -4085
rect 3380 -4165 3410 -4155
rect 3380 -4190 3385 -4165
rect 3405 -4190 3410 -4165
rect 3380 -4230 3410 -4190
rect 3460 -4225 3730 -4220
rect 3900 -4225 3930 -4105
rect 3460 -4230 3930 -4225
rect 3320 -4235 3930 -4230
rect 3320 -4255 3620 -4235
rect 3640 -4255 3930 -4235
rect 3320 -4260 3930 -4255
rect 3278 -4265 3930 -4260
rect 3278 -4280 3460 -4265
rect 3278 -4320 3440 -4280
rect 4100 -4670 4125 -4105
rect 4200 -4130 4225 -4105
rect 4198 -4140 4228 -4130
rect 4198 -4165 4203 -4140
rect 4223 -4165 4228 -4140
rect 4198 -4195 4228 -4165
rect 5075 -4340 5347 -4330
rect 4190 -4350 4230 -4345
rect 4190 -4380 4195 -4350
rect 4225 -4380 4230 -4350
rect 4190 -4385 4230 -4380
rect 4855 -4355 5190 -4340
rect 4855 -4380 4975 -4355
rect 4995 -4360 5190 -4355
rect 5215 -4360 5347 -4340
rect 4995 -4365 5347 -4360
rect 4995 -4380 5105 -4365
rect 4855 -4400 5105 -4380
rect 4100 -4685 4220 -4670
rect 4195 -4725 4220 -4685
rect 4193 -4735 4223 -4725
rect 4193 -4760 4198 -4735
rect 4218 -4760 4223 -4735
rect 4193 -4790 4223 -4760
rect 4185 -4965 4225 -4960
rect 4185 -4995 4190 -4965
rect 4220 -4995 4225 -4965
rect 4185 -5000 4225 -4995
rect 3500 -5100 3780 -5090
rect 3165 -5115 3615 -5100
rect 3165 -5140 3400 -5115
rect 3420 -5120 3615 -5115
rect 3640 -5120 3780 -5100
rect 3420 -5125 3780 -5120
rect 3420 -5140 3530 -5125
rect 3165 -5160 3530 -5140
rect 3165 -5215 3210 -5160
rect 440 -5260 3210 -5215
rect 3745 -5180 3780 -5125
rect 4855 -5180 4885 -4400
rect 5950 -4705 6080 -4690
rect 5950 -4730 5995 -4705
rect 6015 -4720 6340 -4705
rect 6015 -4730 6155 -4720
rect 5950 -4740 6155 -4730
rect 6195 -4740 6340 -4720
rect 5950 -4750 6340 -4740
rect 5950 -5180 5985 -4750
rect 6470 -5065 6515 -3865
rect 7450 -4050 7480 -3405
rect 7550 -3430 7575 -3405
rect 8260 -3395 8265 -3370
rect 8285 -3395 8290 -3370
rect 7548 -3440 7578 -3430
rect 8260 -3435 8290 -3395
rect 9078 -3345 9108 -3335
rect 9078 -3370 9083 -3345
rect 9103 -3370 9108 -3345
rect 9078 -3400 9108 -3370
rect 8340 -3430 8610 -3425
rect 8340 -3435 8800 -3430
rect 7548 -3465 7553 -3440
rect 7573 -3465 7578 -3440
rect 8200 -3440 8800 -3435
rect 8200 -3460 8500 -3440
rect 8520 -3460 8800 -3440
rect 8200 -3465 8800 -3460
rect 7548 -3495 7578 -3465
rect 8158 -3470 8800 -3465
rect 8158 -3485 8340 -3470
rect 8158 -3525 8320 -3485
rect 7540 -3670 7580 -3665
rect 7540 -3700 7545 -3670
rect 7575 -3700 7580 -3670
rect 7540 -3705 7580 -3700
rect 8775 -3865 8800 -3470
rect 9375 -3640 9405 -3630
rect 9375 -3665 9380 -3640
rect 9400 -3665 9405 -3640
rect 9375 -3705 9405 -3665
rect 9685 -3695 9725 -3210
rect 9455 -3705 9725 -3695
rect 9315 -3730 9525 -3705
rect 9575 -3730 9725 -3705
rect 9315 -3735 9725 -3730
rect 9273 -3740 9725 -3735
rect 10755 -3355 10785 -2775
rect 10860 -2800 10885 -2775
rect 10858 -2810 10888 -2800
rect 10858 -2835 10863 -2810
rect 10883 -2835 10888 -2810
rect 10858 -2865 10888 -2835
rect 10850 -3020 10890 -3015
rect 10850 -3050 10855 -3020
rect 10885 -3050 10890 -3020
rect 10850 -3055 10890 -3050
rect 11565 -3145 11595 -2775
rect 11565 -3175 12410 -3145
rect 11565 -3335 11595 -3175
rect 12385 -3300 12410 -3175
rect 10755 -3370 10880 -3355
rect 9273 -3755 9455 -3740
rect 9273 -3795 9435 -3755
rect 10160 -3770 10432 -3760
rect 9775 -3785 10275 -3770
rect 9775 -3810 10060 -3785
rect 10080 -3790 10275 -3785
rect 10300 -3790 10432 -3770
rect 10080 -3795 10432 -3790
rect 10080 -3810 10190 -3795
rect 9775 -3830 10190 -3810
rect 8775 -3890 9100 -3865
rect 9075 -3930 9100 -3890
rect 9073 -3940 9103 -3930
rect 9073 -3965 9078 -3940
rect 9098 -3965 9103 -3940
rect 9073 -3995 9103 -3965
rect 7205 -4070 7530 -4050
rect 6685 -4130 6715 -4120
rect 6685 -4155 6690 -4130
rect 6710 -4155 6715 -4130
rect 6685 -4195 6715 -4155
rect 6765 -4190 7035 -4185
rect 7205 -4190 7235 -4070
rect 6765 -4195 7235 -4190
rect 6625 -4200 7235 -4195
rect 6625 -4220 6925 -4200
rect 6945 -4220 7235 -4200
rect 6625 -4225 7235 -4220
rect 6583 -4230 7235 -4225
rect 6583 -4245 6765 -4230
rect 6583 -4285 6745 -4245
rect 7410 -4625 7440 -4070
rect 7505 -4095 7530 -4070
rect 7503 -4105 7533 -4095
rect 7503 -4130 7508 -4105
rect 7528 -4130 7533 -4105
rect 7503 -4160 7533 -4130
rect 8380 -4305 8652 -4295
rect 7495 -4315 7535 -4310
rect 7495 -4345 7500 -4315
rect 7530 -4345 7535 -4315
rect 7495 -4350 7535 -4345
rect 8160 -4320 8495 -4305
rect 8160 -4345 8280 -4320
rect 8300 -4325 8495 -4320
rect 8520 -4325 8652 -4305
rect 8300 -4330 8652 -4325
rect 8300 -4345 8410 -4330
rect 8160 -4365 8410 -4345
rect 7410 -4650 7525 -4625
rect 7500 -4690 7525 -4650
rect 7498 -4700 7528 -4690
rect 7498 -4725 7503 -4700
rect 7523 -4725 7528 -4700
rect 7498 -4755 7528 -4725
rect 7490 -4930 7530 -4925
rect 7490 -4960 7495 -4930
rect 7525 -4960 7530 -4930
rect 7490 -4965 7530 -4960
rect 6805 -5065 7085 -5055
rect 6470 -5080 6920 -5065
rect 6470 -5105 6705 -5080
rect 6725 -5085 6920 -5080
rect 6945 -5085 7085 -5065
rect 6725 -5090 7085 -5085
rect 6725 -5105 6835 -5090
rect 6470 -5125 6835 -5105
rect 6470 -5180 6515 -5125
rect 3745 -5225 6515 -5180
rect 7050 -5145 7085 -5090
rect 8160 -5145 8190 -4365
rect 9265 -4670 9395 -4655
rect 9265 -4695 9310 -4670
rect 9330 -4685 9655 -4670
rect 9330 -4695 9470 -4685
rect 9265 -4705 9470 -4695
rect 9510 -4705 9655 -4685
rect 9265 -4715 9655 -4705
rect 9365 -5145 9400 -4715
rect 9775 -5030 9820 -3830
rect 10755 -4015 10785 -3370
rect 10855 -3395 10880 -3370
rect 11565 -3360 11570 -3335
rect 11590 -3360 11595 -3335
rect 10853 -3405 10883 -3395
rect 11565 -3400 11595 -3360
rect 12383 -3310 12413 -3300
rect 12383 -3335 12388 -3310
rect 12408 -3335 12413 -3310
rect 12383 -3365 12413 -3335
rect 11645 -3395 11915 -3390
rect 11645 -3400 12105 -3395
rect 10853 -3430 10858 -3405
rect 10878 -3430 10883 -3405
rect 11505 -3405 12105 -3400
rect 11505 -3425 11805 -3405
rect 11825 -3425 12105 -3405
rect 11505 -3430 12105 -3425
rect 10853 -3460 10883 -3430
rect 11463 -3435 12105 -3430
rect 11463 -3450 11645 -3435
rect 11463 -3490 11625 -3450
rect 10845 -3635 10885 -3630
rect 10845 -3665 10850 -3635
rect 10880 -3665 10885 -3635
rect 10845 -3670 10885 -3665
rect 12080 -3830 12105 -3435
rect 12080 -3855 12405 -3830
rect 12380 -3895 12405 -3855
rect 12378 -3905 12408 -3895
rect 12378 -3930 12383 -3905
rect 12403 -3930 12408 -3905
rect 12378 -3960 12408 -3930
rect 10510 -4035 10835 -4015
rect 9990 -4095 10020 -4085
rect 9990 -4120 9995 -4095
rect 10015 -4120 10020 -4095
rect 9990 -4160 10020 -4120
rect 10070 -4155 10340 -4150
rect 10510 -4155 10540 -4035
rect 10070 -4160 10540 -4155
rect 9930 -4165 10540 -4160
rect 9930 -4185 10230 -4165
rect 10250 -4185 10540 -4165
rect 9930 -4190 10540 -4185
rect 9888 -4195 10540 -4190
rect 9888 -4210 10070 -4195
rect 9888 -4250 10050 -4210
rect 10715 -4590 10755 -4035
rect 10810 -4060 10835 -4035
rect 10808 -4070 10838 -4060
rect 10808 -4095 10813 -4070
rect 10833 -4095 10838 -4070
rect 10808 -4125 10838 -4095
rect 12885 -4120 12955 -2615
rect 13215 -3105 13245 -1755
rect 13215 -3130 13220 -3105
rect 13240 -3130 13245 -3105
rect 13645 -3065 13675 -3005
rect 13645 -3090 13650 -3065
rect 13670 -3090 13675 -3065
rect 13645 -3130 13675 -3090
rect 13725 -3130 13985 -3120
rect 13215 -3170 13245 -3130
rect 13585 -3155 13795 -3130
rect 13845 -3155 13985 -3130
rect 13585 -3160 13985 -3155
rect 13295 -3165 13985 -3160
rect 13295 -3170 13725 -3165
rect 13155 -3195 13365 -3170
rect 13415 -3180 13725 -3170
rect 13415 -3195 13705 -3180
rect 13155 -3200 13705 -3195
rect 13113 -3205 13705 -3200
rect 13113 -3220 13295 -3205
rect 13543 -3220 13705 -3205
rect 13113 -3260 13275 -3220
rect 13525 -4095 13665 -4080
rect 13525 -4120 13580 -4095
rect 13600 -4110 13925 -4095
rect 13600 -4120 13740 -4110
rect 12885 -4135 13235 -4120
rect 13525 -4130 13740 -4120
rect 13780 -4130 13925 -4110
rect 13525 -4135 13925 -4130
rect 12885 -4160 13150 -4135
rect 13170 -4140 13925 -4135
rect 13170 -4150 13555 -4140
rect 13170 -4160 13310 -4150
rect 12885 -4170 13310 -4160
rect 13350 -4170 13555 -4150
rect 12885 -4175 13555 -4170
rect 11685 -4270 11957 -4260
rect 10800 -4280 10840 -4275
rect 10800 -4310 10805 -4280
rect 10835 -4310 10840 -4280
rect 10800 -4315 10840 -4310
rect 11465 -4285 11800 -4270
rect 11465 -4310 11585 -4285
rect 11605 -4290 11800 -4285
rect 11825 -4290 11957 -4270
rect 11605 -4295 11957 -4290
rect 11605 -4310 11715 -4295
rect 11465 -4330 11715 -4310
rect 10715 -4615 10830 -4590
rect 10805 -4655 10830 -4615
rect 10803 -4665 10833 -4655
rect 10803 -4690 10808 -4665
rect 10828 -4690 10833 -4665
rect 10803 -4720 10833 -4690
rect 10795 -4895 10835 -4890
rect 10795 -4925 10800 -4895
rect 10830 -4925 10835 -4895
rect 10795 -4930 10835 -4925
rect 10110 -5030 10390 -5020
rect 9775 -5045 10225 -5030
rect 9775 -5070 10010 -5045
rect 10030 -5050 10225 -5045
rect 10250 -5050 10390 -5030
rect 10030 -5055 10390 -5050
rect 10030 -5070 10140 -5055
rect 9775 -5090 10140 -5070
rect 9775 -5145 9820 -5090
rect 7050 -5190 9820 -5145
rect 10355 -5110 10390 -5055
rect 11465 -5110 11495 -4330
rect 12885 -5110 12955 -4175
rect 13105 -4180 13555 -4175
rect 10355 -5155 12955 -5110
rect 5950 -5230 5985 -5225
rect 9355 -5305 9385 -5295
rect 9355 -5330 9360 -5305
rect 9380 -5330 9385 -5305
rect 9355 -5370 9385 -5330
rect 9435 -5370 9695 -5360
rect 9295 -5395 9505 -5370
rect 9555 -5395 9695 -5370
rect 9295 -5400 9695 -5395
rect 9253 -5405 9695 -5400
rect 6250 -5425 6280 -5415
rect 6250 -5450 6255 -5425
rect 6275 -5450 6280 -5425
rect 6250 -5490 6280 -5450
rect 9253 -5420 9435 -5405
rect 9253 -5460 9415 -5420
rect 6585 -5480 9375 -5460
rect 6330 -5490 9375 -5480
rect 6190 -5515 6400 -5490
rect 6450 -5515 9375 -5490
rect 6190 -5520 9375 -5515
rect 2805 -5530 2835 -5520
rect 2805 -5555 2810 -5530
rect 2830 -5555 2835 -5530
rect 2805 -5595 2835 -5555
rect 6148 -5525 9375 -5520
rect 6148 -5540 6330 -5525
rect 6148 -5580 6310 -5540
rect 3140 -5585 6230 -5580
rect 2885 -5595 6230 -5585
rect 2745 -5620 2955 -5595
rect 3005 -5620 6230 -5595
rect 2745 -5625 6230 -5620
rect -370 -5630 -160 -5625
rect 2703 -5630 6230 -5625
rect -370 -5645 2885 -5630
rect -370 -5680 2865 -5645
rect 2703 -5685 2865 -5680
rect 9245 -6335 9375 -6320
rect 10480 -6330 10545 -5155
rect 9995 -6335 10545 -6330
rect 9245 -6360 9290 -6335
rect 9310 -6350 10545 -6335
rect 9310 -6360 9450 -6350
rect 9245 -6370 9450 -6360
rect 9490 -6370 10545 -6350
rect 9245 -6380 10545 -6370
rect 6140 -6455 6270 -6440
rect 9550 -6455 9580 -6380
rect 6140 -6480 6185 -6455
rect 6205 -6470 9580 -6455
rect 6205 -6480 6345 -6470
rect 6140 -6490 6345 -6480
rect 6385 -6490 9580 -6470
rect 6140 -6500 9580 -6490
rect 2695 -6560 2825 -6545
rect 6140 -6560 6200 -6500
rect 2695 -6585 2740 -6560
rect 2760 -6575 6200 -6560
rect 2760 -6585 2900 -6575
rect 2695 -6595 2900 -6585
rect 2940 -6595 6200 -6575
rect 2695 -6605 6200 -6595
<< via1 >>
rect 360 -2360 390 -2355
rect 360 -2380 365 -2360
rect 365 -2380 385 -2360
rect 385 -2380 390 -2360
rect 360 -2385 390 -2380
rect 1850 -2370 1880 -2365
rect 1850 -2390 1855 -2370
rect 1855 -2390 1875 -2370
rect 1875 -2390 1880 -2370
rect 1850 -2395 1880 -2390
rect 2980 -2340 3010 -2335
rect 2980 -2360 2985 -2340
rect 2985 -2360 3005 -2340
rect 3005 -2360 3010 -2340
rect 2980 -2365 3010 -2360
rect 3665 -2325 3695 -2320
rect 3665 -2345 3670 -2325
rect 3670 -2345 3690 -2325
rect 3690 -2345 3695 -2325
rect 3665 -2350 3695 -2345
rect 5155 -2335 5185 -2330
rect 5155 -2355 5160 -2335
rect 5160 -2355 5180 -2335
rect 5180 -2355 5185 -2335
rect 5155 -2360 5185 -2355
rect 6285 -2305 6315 -2300
rect 6285 -2325 6290 -2305
rect 6290 -2325 6310 -2305
rect 6310 -2325 6315 -2305
rect 6285 -2330 6315 -2325
rect 6970 -2290 7000 -2285
rect 6970 -2310 6975 -2290
rect 6975 -2310 6995 -2290
rect 6995 -2310 7000 -2290
rect 6970 -2315 7000 -2310
rect 8460 -2300 8490 -2295
rect 8460 -2320 8465 -2300
rect 8465 -2320 8485 -2300
rect 8485 -2320 8490 -2300
rect 8460 -2325 8490 -2320
rect 9590 -2270 9620 -2265
rect 9590 -2290 9595 -2270
rect 9595 -2290 9615 -2270
rect 9615 -2290 9620 -2270
rect 9590 -2295 9620 -2290
rect 10275 -2255 10305 -2250
rect 10275 -2275 10280 -2255
rect 10280 -2275 10300 -2255
rect 10300 -2275 10305 -2255
rect 10275 -2280 10305 -2275
rect 11765 -2265 11795 -2260
rect 11765 -2285 11770 -2265
rect 11770 -2285 11790 -2265
rect 11790 -2285 11795 -2265
rect 11765 -2290 11795 -2285
rect 12895 -2235 12925 -2230
rect 12895 -2255 12900 -2235
rect 12900 -2255 12920 -2235
rect 12920 -2255 12925 -2235
rect 12895 -2260 12925 -2255
rect 830 -2455 860 -2450
rect 830 -2475 835 -2455
rect 835 -2475 855 -2455
rect 855 -2475 860 -2455
rect 830 -2480 860 -2475
rect 4135 -2420 4165 -2415
rect 4135 -2440 4140 -2420
rect 4140 -2440 4160 -2420
rect 4160 -2440 4165 -2420
rect 4135 -2445 4165 -2440
rect 7440 -2385 7470 -2380
rect 7440 -2405 7445 -2385
rect 7445 -2405 7465 -2385
rect 7465 -2405 7470 -2385
rect 7440 -2410 7470 -2405
rect 10745 -2350 10775 -2345
rect 10745 -2370 10750 -2350
rect 10750 -2370 10770 -2350
rect 10770 -2370 10775 -2350
rect 10745 -2375 10775 -2370
rect 940 -3130 970 -3125
rect 940 -3150 945 -3130
rect 945 -3150 965 -3130
rect 965 -3150 970 -3130
rect 940 -3155 970 -3150
rect 935 -3745 965 -3740
rect 935 -3765 940 -3745
rect 940 -3765 960 -3745
rect 960 -3765 965 -3745
rect 935 -3770 965 -3765
rect 4245 -3095 4275 -3090
rect 4245 -3115 4250 -3095
rect 4250 -3115 4270 -3095
rect 4270 -3115 4275 -3095
rect 4245 -3120 4275 -3115
rect 890 -4390 920 -4385
rect 890 -4410 895 -4390
rect 895 -4410 915 -4390
rect 915 -4410 920 -4390
rect 890 -4415 920 -4410
rect 885 -5005 915 -5000
rect 885 -5025 890 -5005
rect 890 -5025 910 -5005
rect 910 -5025 915 -5005
rect 885 -5030 915 -5025
rect 4240 -3710 4270 -3705
rect 4240 -3730 4245 -3710
rect 4245 -3730 4265 -3710
rect 4265 -3730 4270 -3710
rect 4240 -3735 4270 -3730
rect 7550 -3060 7580 -3055
rect 7550 -3080 7555 -3060
rect 7555 -3080 7575 -3060
rect 7575 -3080 7580 -3060
rect 7550 -3085 7580 -3080
rect 4195 -4355 4225 -4350
rect 4195 -4375 4200 -4355
rect 4200 -4375 4220 -4355
rect 4220 -4375 4225 -4355
rect 4195 -4380 4225 -4375
rect 4190 -4970 4220 -4965
rect 4190 -4990 4195 -4970
rect 4195 -4990 4215 -4970
rect 4215 -4990 4220 -4970
rect 4190 -4995 4220 -4990
rect 7545 -3675 7575 -3670
rect 7545 -3695 7550 -3675
rect 7550 -3695 7570 -3675
rect 7570 -3695 7575 -3675
rect 7545 -3700 7575 -3695
rect 10855 -3025 10885 -3020
rect 10855 -3045 10860 -3025
rect 10860 -3045 10880 -3025
rect 10880 -3045 10885 -3025
rect 10855 -3050 10885 -3045
rect 7500 -4320 7530 -4315
rect 7500 -4340 7505 -4320
rect 7505 -4340 7525 -4320
rect 7525 -4340 7530 -4320
rect 7500 -4345 7530 -4340
rect 7495 -4935 7525 -4930
rect 7495 -4955 7500 -4935
rect 7500 -4955 7520 -4935
rect 7520 -4955 7525 -4935
rect 7495 -4960 7525 -4955
rect 10850 -3640 10880 -3635
rect 10850 -3660 10855 -3640
rect 10855 -3660 10875 -3640
rect 10875 -3660 10880 -3640
rect 10850 -3665 10880 -3660
rect 10805 -4285 10835 -4280
rect 10805 -4305 10810 -4285
rect 10810 -4305 10830 -4285
rect 10830 -4305 10835 -4285
rect 10805 -4310 10835 -4305
rect 10800 -4900 10830 -4895
rect 10800 -4920 10805 -4900
rect 10805 -4920 10825 -4900
rect 10825 -4920 10830 -4900
rect 10800 -4925 10830 -4920
<< metal2 >>
rect 12890 -2230 12930 -2225
rect 10270 -2250 10310 -2245
rect 9585 -2265 9625 -2260
rect 6965 -2285 7005 -2280
rect 6280 -2300 6320 -2295
rect 3660 -2320 3700 -2315
rect 2975 -2335 3015 -2330
rect 355 -2355 395 -2350
rect 355 -2385 360 -2355
rect 390 -2385 395 -2355
rect 355 -2390 395 -2385
rect 1845 -2365 1885 -2360
rect 355 -2825 385 -2390
rect 1845 -2395 1850 -2365
rect 1880 -2370 1885 -2365
rect 2975 -2365 2980 -2335
rect 3010 -2365 3135 -2335
rect 2975 -2370 3015 -2365
rect 1880 -2390 2020 -2370
rect 1880 -2395 1885 -2390
rect 1845 -2400 1885 -2395
rect 825 -2450 865 -2445
rect 825 -2480 830 -2450
rect 860 -2480 865 -2450
rect 825 -2485 865 -2480
rect 845 -2790 865 -2485
rect 1995 -2790 2020 -2390
rect 845 -2805 1140 -2790
rect 355 -2845 570 -2825
rect 550 -3130 570 -2845
rect 935 -3125 975 -3120
rect 935 -3130 940 -3125
rect 550 -3150 940 -3130
rect 935 -3155 940 -3150
rect 970 -3155 975 -3125
rect 935 -3160 975 -3155
rect 930 -3740 970 -3735
rect 930 -3770 935 -3740
rect 965 -3745 970 -3740
rect 1120 -3745 1140 -2805
rect 965 -3765 1140 -3745
rect 1230 -2820 2020 -2790
rect 965 -3770 970 -3765
rect 930 -3775 970 -3770
rect 885 -4385 925 -4380
rect 885 -4415 890 -4385
rect 920 -4390 925 -4385
rect 1230 -4390 1250 -2820
rect 3100 -2880 3135 -2365
rect 3660 -2350 3665 -2320
rect 3695 -2350 3700 -2320
rect 3660 -2355 3700 -2350
rect 5150 -2330 5190 -2325
rect 3660 -2790 3690 -2355
rect 5150 -2360 5155 -2330
rect 5185 -2335 5190 -2330
rect 6280 -2330 6285 -2300
rect 6315 -2330 6440 -2300
rect 6280 -2335 6320 -2330
rect 5185 -2355 5325 -2335
rect 5185 -2360 5190 -2355
rect 5150 -2365 5190 -2360
rect 4130 -2415 4170 -2410
rect 4130 -2445 4135 -2415
rect 4165 -2445 4170 -2415
rect 4130 -2450 4170 -2445
rect 4150 -2755 4170 -2450
rect 5300 -2755 5325 -2355
rect 4150 -2770 4445 -2755
rect 3660 -2810 3875 -2790
rect 920 -4415 1250 -4390
rect 1390 -2910 3135 -2880
rect 885 -4420 925 -4415
rect 880 -5000 920 -4995
rect 1390 -5000 1410 -2910
rect 3855 -3095 3875 -2810
rect 4240 -3090 4280 -3085
rect 4240 -3095 4245 -3090
rect 3855 -3115 4245 -3095
rect 4240 -3120 4245 -3115
rect 4275 -3120 4280 -3090
rect 4240 -3125 4280 -3120
rect 4235 -3705 4275 -3700
rect 4235 -3735 4240 -3705
rect 4270 -3710 4275 -3705
rect 4425 -3710 4445 -2770
rect 4270 -3730 4445 -3710
rect 4535 -2785 5325 -2755
rect 4270 -3735 4275 -3730
rect 4235 -3740 4275 -3735
rect 4190 -4350 4230 -4345
rect 4190 -4380 4195 -4350
rect 4225 -4355 4230 -4350
rect 4535 -4355 4555 -2785
rect 6405 -2845 6440 -2330
rect 6965 -2315 6970 -2285
rect 7000 -2315 7005 -2285
rect 6965 -2320 7005 -2315
rect 8455 -2295 8495 -2290
rect 6965 -2755 6995 -2320
rect 8455 -2325 8460 -2295
rect 8490 -2300 8495 -2295
rect 9585 -2295 9590 -2265
rect 9620 -2295 9745 -2265
rect 9585 -2300 9625 -2295
rect 8490 -2320 8630 -2300
rect 8490 -2325 8495 -2320
rect 8455 -2330 8495 -2325
rect 7435 -2380 7475 -2375
rect 7435 -2410 7440 -2380
rect 7470 -2410 7475 -2380
rect 7435 -2415 7475 -2410
rect 7455 -2720 7475 -2415
rect 8605 -2720 8630 -2320
rect 7455 -2735 7750 -2720
rect 6965 -2775 7180 -2755
rect 4225 -4380 4555 -4355
rect 4695 -2875 6440 -2845
rect 4190 -4385 4230 -4380
rect 4185 -4965 4225 -4960
rect 4695 -4965 4715 -2875
rect 7160 -3060 7180 -2775
rect 7545 -3055 7585 -3050
rect 7545 -3060 7550 -3055
rect 7160 -3080 7550 -3060
rect 7545 -3085 7550 -3080
rect 7580 -3085 7585 -3055
rect 7545 -3090 7585 -3085
rect 7540 -3670 7580 -3665
rect 7540 -3700 7545 -3670
rect 7575 -3675 7580 -3670
rect 7730 -3675 7750 -2735
rect 7575 -3695 7750 -3675
rect 7840 -2750 8630 -2720
rect 7575 -3700 7580 -3695
rect 7540 -3705 7580 -3700
rect 7495 -4315 7535 -4310
rect 7495 -4345 7500 -4315
rect 7530 -4320 7535 -4315
rect 7840 -4320 7860 -2750
rect 9710 -2810 9745 -2295
rect 10270 -2280 10275 -2250
rect 10305 -2280 10310 -2250
rect 10270 -2285 10310 -2280
rect 11760 -2260 11800 -2255
rect 10270 -2720 10300 -2285
rect 11760 -2290 11765 -2260
rect 11795 -2265 11800 -2260
rect 12890 -2260 12895 -2230
rect 12925 -2260 13050 -2230
rect 12890 -2265 12930 -2260
rect 11795 -2285 11935 -2265
rect 11795 -2290 11800 -2285
rect 11760 -2295 11800 -2290
rect 10740 -2345 10780 -2340
rect 10740 -2375 10745 -2345
rect 10775 -2375 10780 -2345
rect 10740 -2380 10780 -2375
rect 10760 -2685 10780 -2380
rect 11910 -2685 11935 -2285
rect 10760 -2700 11055 -2685
rect 10270 -2740 10485 -2720
rect 7530 -4345 7860 -4320
rect 8000 -2840 9745 -2810
rect 7495 -4350 7535 -4345
rect 7490 -4930 7530 -4925
rect 8000 -4930 8020 -2840
rect 10465 -3025 10485 -2740
rect 10850 -3020 10890 -3015
rect 10850 -3025 10855 -3020
rect 10465 -3045 10855 -3025
rect 10850 -3050 10855 -3045
rect 10885 -3050 10890 -3020
rect 10850 -3055 10890 -3050
rect 10845 -3635 10885 -3630
rect 10845 -3665 10850 -3635
rect 10880 -3640 10885 -3635
rect 11035 -3640 11055 -2700
rect 10880 -3660 11055 -3640
rect 11145 -2715 11935 -2685
rect 10880 -3665 10885 -3660
rect 10845 -3670 10885 -3665
rect 10800 -4280 10840 -4275
rect 10800 -4310 10805 -4280
rect 10835 -4285 10840 -4280
rect 11145 -4285 11165 -2715
rect 13015 -2775 13050 -2260
rect 10835 -4310 11165 -4285
rect 11305 -2805 13050 -2775
rect 10800 -4315 10840 -4310
rect 10795 -4895 10835 -4890
rect 11305 -4895 11325 -2805
rect 10795 -4925 10800 -4895
rect 10830 -4920 11325 -4895
rect 10830 -4925 10835 -4920
rect 10795 -4930 10835 -4925
rect 7490 -4960 7495 -4930
rect 7525 -4955 8020 -4930
rect 7525 -4960 7530 -4955
rect 7490 -4965 7530 -4960
rect 4185 -4995 4190 -4965
rect 4220 -4990 4715 -4965
rect 4220 -4995 4225 -4990
rect 4185 -5000 4225 -4995
rect 880 -5030 885 -5000
rect 915 -5025 1410 -5000
rect 915 -5030 920 -5025
rect 880 -5035 920 -5030
<< labels >>
rlabel viali 195 -1885 240 -1860 1 Vdd
rlabel viali 185 -2755 235 -2730 1 gnd
rlabel metal1 610 -1910 770 -1855 1 Vdd
rlabel metal1 610 -2755 810 -2700 1 gnd
rlabel metal1 1780 -2750 1840 -2720 1 gnd
rlabel metal1 1780 -1885 1840 -1855 1 Vdd
rlabel locali 1835 -2415 1890 -2340 1 AND0
rlabel locali 1495 -2400 1575 -2360 1 net10
rlabel locali 2560 -2370 2640 -2330 1 net1
rlabel locali 2965 -2370 3020 -2325 1 OR0
rlabel metal1 2195 -2755 2395 -2700 1 gnd
rlabel metal1 2195 -1910 2355 -1855 1 Vdd
rlabel metal1 2910 -2720 2970 -2690 1 gnd
rlabel metal1 2910 -1855 2970 -1825 1 Vdd
rlabel metal1 345 -3900 405 -3870 1 gnd
rlabel metal1 345 -3035 405 -3005 1 Vdd
rlabel metal1 295 -5160 355 -5130 1 gnd
rlabel metal1 295 -4295 355 -4265 1 Vdd
rlabel metal1 1870 -3535 1930 -3505 1 Vdd
rlabel metal1 1870 -4400 1930 -4370 1 gnd
rlabel metal2 355 -2390 395 -2350 1 NAND0
rlabel metal2 825 -2485 865 -2445 1 NOR0
rlabel poly 1815 -4055 1890 -4005 1 S1_0
rlabel ndiff 1280 -2630 1330 -2515 1 net9
rlabel ndiff 195 -2620 245 -2505 1 net21
rlabel pdiff 2270 -2260 2325 -2030 1 net2
rlabel viali 3500 -1850 3545 -1825 1 Vdd
rlabel viali 3490 -2720 3540 -2695 1 gnd
rlabel metal1 3915 -1875 4075 -1820 1 Vdd
rlabel metal1 3915 -2720 4115 -2665 1 gnd
rlabel metal1 5085 -2715 5145 -2685 1 gnd
rlabel metal1 5085 -1850 5145 -1820 1 Vdd
rlabel metal1 5500 -2720 5700 -2665 1 gnd
rlabel metal1 5500 -1875 5660 -1820 1 Vdd
rlabel metal1 6215 -2685 6275 -2655 1 gnd
rlabel metal1 6215 -1820 6275 -1790 1 Vdd
rlabel metal1 3650 -3865 3710 -3835 1 gnd
rlabel metal1 3650 -3000 3710 -2970 1 Vdd
rlabel metal1 3600 -5125 3660 -5095 1 gnd
rlabel metal1 3600 -4260 3660 -4230 1 Vdd
rlabel metal1 5175 -3500 5235 -3470 1 Vdd
rlabel metal1 5175 -4365 5235 -4335 1 gnd
rlabel viali 6805 -1815 6850 -1790 1 Vdd
rlabel viali 6795 -2685 6845 -2660 1 gnd
rlabel metal1 7220 -1840 7380 -1785 1 Vdd
rlabel metal1 7220 -2685 7420 -2630 1 gnd
rlabel metal1 8390 -2680 8450 -2650 1 gnd
rlabel metal1 8390 -1815 8450 -1785 1 Vdd
rlabel metal1 8805 -2685 9005 -2630 1 gnd
rlabel metal1 8805 -1840 8965 -1785 1 Vdd
rlabel metal1 9520 -2650 9580 -2620 1 gnd
rlabel metal1 9520 -1785 9580 -1755 1 Vdd
rlabel metal1 6955 -3830 7015 -3800 1 gnd
rlabel metal1 6955 -2965 7015 -2935 1 Vdd
rlabel metal1 6905 -5090 6965 -5060 1 gnd
rlabel metal1 6905 -4225 6965 -4195 1 Vdd
rlabel metal1 8480 -3465 8540 -3435 1 Vdd
rlabel metal1 8480 -4330 8540 -4300 1 gnd
rlabel metal1 11785 -4295 11845 -4265 1 gnd
rlabel metal1 11785 -3430 11845 -3400 1 Vdd
rlabel metal1 10210 -4190 10270 -4160 1 Vdd
rlabel metal1 10210 -5055 10270 -5025 1 gnd
rlabel metal1 10260 -2930 10320 -2900 1 Vdd
rlabel metal1 10260 -3795 10320 -3765 1 gnd
rlabel metal1 12825 -1750 12885 -1720 1 Vdd
rlabel metal1 12825 -2615 12885 -2585 1 gnd
rlabel metal1 12110 -1805 12270 -1750 1 Vdd
rlabel metal1 12110 -2650 12310 -2595 1 gnd
rlabel metal1 11695 -1780 11755 -1750 1 Vdd
rlabel metal1 11695 -2645 11755 -2615 1 gnd
rlabel metal1 10525 -2650 10725 -2595 1 gnd
rlabel metal1 10525 -1805 10685 -1750 1 Vdd
rlabel viali 10100 -2650 10150 -2625 1 gnd
rlabel viali 10110 -1780 10155 -1755 1 Vdd
rlabel metal1 120 -2255 170 -2210 1 A0_0
rlabel metal1 210 -2415 250 -2375 1 B0_0
rlabel pdiff 690 -2255 745 -2025 1 net17
rlabel metal1 620 -2415 660 -2385 1 A0_1
rlabel metal1 710 -2495 750 -2465 1 B0_1
rlabel metal1 1205 -2265 1255 -2220 1 A0_2
rlabel poly 1295 -2425 1345 -2380 1 B0_2
rlabel metal1 2205 -2415 2245 -2385 1 A0_3
rlabel metal1 2295 -2495 2335 -2465 1 B0_3
rlabel metal1 3425 -2220 3475 -2175 1 A1_0
rlabel poly 3515 -2380 3565 -2335 1 B1_0
rlabel metal2 3660 -2355 3700 -2315 1 NAND1
rlabel ndiff 3500 -2585 3550 -2470 1 net22
rlabel metal2 4130 -2450 4170 -2410 1 NOR1
rlabel pdiff 3995 -2220 4050 -1990 1 net18
rlabel metal1 3925 -2380 3965 -2350 1 A1_1
rlabel metal1 4015 -2460 4055 -2430 1 B1_1
rlabel metal1 4510 -2230 4560 -2185 1 A1_2
rlabel poly 4600 -2390 4650 -2345 1 B1_2
rlabel locali 4795 -2365 4905 -2325 1 net12
rlabel ndiff 4585 -2595 4635 -2480 1 net11
rlabel locali 5140 -2380 5195 -2305 1 AND1
rlabel pdiff 5575 -2225 5630 -1995 1 net4
rlabel locali 5865 -2335 5945 -2295 1 net3
rlabel locali 6270 -2335 6325 -2290 1 OR1
rlabel metal2 6965 -2320 7005 -2280 1 NAN2
rlabel metal1 6730 -2185 6780 -2140 1 A2_0
rlabel poly 6820 -2345 6870 -2300 1 B2_0
rlabel ndiff 6805 -2550 6855 -2435 1 net23
rlabel metal2 7435 -2415 7475 -2375 1 NOR2
rlabel metal1 7230 -2345 7270 -2315 1 A2_1
rlabel metal1 7320 -2425 7360 -2395 1 B2_1
rlabel pdiff 7300 -2185 7355 -1955 1 net19
rlabel locali 8445 -2345 8500 -2270 1 AND2
rlabel ndiff 7890 -2560 7940 -2445 1 net13
rlabel metal1 7815 -2195 7865 -2150 1 A2_2
rlabel poly 7905 -2355 7955 -2310 1 B2_2
rlabel locali 8105 -2330 8185 -2290 1 net14
rlabel locali 9575 -2300 9630 -2255 1 OR2
rlabel locali 9170 -2300 9250 -2260 1 net5
rlabel metal1 8815 -2345 8855 -2315 1 A2_3
rlabel metal1 8905 -2425 8945 -2395 1 B2_3
rlabel pdiff 8880 -2190 8935 -1960 1 net6
rlabel ndiff 10110 -2515 10160 -2400 1 net24
rlabel poly 10125 -2310 10175 -2265 1 B3_0
rlabel metal1 10035 -2150 10085 -2105 1 A3_0
rlabel metal2 10270 -2285 10310 -2245 1 NAND3
rlabel metal1 10535 -2310 10575 -2280 1 A3_1
rlabel metal1 10625 -2390 10665 -2360 1 B3_1
rlabel pdiff 10605 -2150 10660 -1920 1 net20
rlabel metal2 10740 -2380 10780 -2340 1 NOR3
rlabel locali 11750 -2310 11805 -2235 1 AND3
rlabel locali 11410 -2295 11490 -2255 1 net16
rlabel ndiff 11195 -2525 11245 -2410 1 net15
rlabel metal1 11120 -2160 11170 -2115 1 A3_2
rlabel poly 11210 -2320 11260 -2275 1 B3_2
rlabel metal1 12120 -2310 12160 -2280 1 A3_3
rlabel metal1 12210 -2390 12250 -2360 1 B3_3
rlabel pdiff 12185 -2155 12240 -1925 1 net8
rlabel locali 12475 -2265 12555 -2225 1 net7
rlabel locali 12880 -2265 12935 -2220 1 OR3
rlabel poly 290 -3555 365 -3505 1 S0_0
rlabel locali 540 -3585 585 -3565 1 net46
rlabel locali 1035 -3415 1105 -3375 1 net47
rlabel locali 435 -4845 490 -4825 1 net52
rlabel poly 240 -4815 315 -4765 1 S0_1
rlabel locali 1005 -4675 1090 -4630 1 net50
rlabel locali 2025 -4085 2075 -4065 1 net49
rlabel locali 2585 -3915 2635 -3875 1 net48
rlabel poly 3595 -3520 3670 -3470 1 S0_2
rlabel poly 3545 -4780 3620 -4730 1 S0_3
rlabel locali 3800 -3550 3860 -3530 1 net39
rlabel locali 4375 -4640 4445 -4600 1 net43
rlabel locali 4340 -3380 4410 -3340 1 net40
rlabel poly 5120 -4020 5195 -3970 1 S1_1
rlabel locali 5300 -4050 5375 -4030 1 net42
rlabel locali 5890 -3880 5940 -3840 1 net41
rlabel poly 6900 -3485 6975 -3435 1 S0_4
rlabel poly 6850 -4745 6925 -4695 1 S0_5
rlabel locali 7090 -3515 7125 -3495 1 net32
rlabel locali 7025 -4775 7105 -4755 1 net38
rlabel locali 7645 -3345 7695 -3305 1 net33
rlabel locali 7600 -4605 7710 -4565 1 net36
rlabel locali 8540 -4020 8590 -3990 1 net35
rlabel poly 8425 -3985 8500 -3935 1 S1_2
rlabel locali 9195 -3845 9245 -3805 1 net34
rlabel poly 10205 -3450 10280 -3400 1 S0_6
rlabel poly 10155 -4710 10230 -4660 1 S0_7
rlabel locali 10320 -3480 10360 -3440 1 net25
rlabel locali 10265 -4745 10315 -4705 1 net31
rlabel locali 10955 -3310 11000 -3270 1 net26
rlabel locali 10920 -4570 10980 -4535 1 net29
rlabel poly 11730 -3950 11805 -3900 1 S1_3
rlabel locali 11840 -3985 11890 -3945 1 net28
rlabel locali 12500 -3810 12550 -3770 1 net27
rlabel locali 3735 -4810 3785 -4790 1 net45
rlabel locali 13845 -3785 13920 -3740 1 F3
rlabel locali 13540 -3780 13630 -3740 1 net30
rlabel locali 9585 -4375 9635 -4315 1 net37
rlabel locali 6275 -4385 6320 -4325 1 net44
rlabel locali 2940 -4425 2995 -4370 1 net51
rlabel locali 3010 -6255 3080 -6185 1 F0
rlabel locali 6460 -6145 6515 -6080 1 F1
rlabel locali 9565 -6030 9630 -5955 1 F2
rlabel viali 2880 -3800 2930 -3775 1 Vdd
rlabel viali 2955 -5620 3005 -5595 1 Vdd
rlabel metal1 6400 -5520 6450 -5490 1 Vdd
rlabel metal1 9505 -5395 9555 -5365 1 Vdd
rlabel metal1 13365 -3195 13415 -3165 1 Vdd
rlabel metal1 13800 -3155 13850 -3125 1 Vdd
rlabel viali 11195 -1790 11240 -1765 1 Vdd
rlabel viali 6210 -3765 6260 -3740 1 Vdd
rlabel viali 9525 -3730 9575 -3705 1 Vdd
rlabel viali 1280 -1895 1325 -1870 1 Vdd
rlabel nwell 2690 -1785 2720 -1750 1 Vdd
rlabel metal1 5510 -2380 5550 -2350 1 A1_3
rlabel metal1 5600 -2460 5640 -2430 1 B1_3
<< end >>
